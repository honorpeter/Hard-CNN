`timescale 1ns / 1ps
// convolution layer control module

module conv_ctrl#(parameter WIDTH = 9)
(
    input clk,
    input rst_n,
    // data
    input [WIDTH-1:0] data_in [31:0],

    output
);

initial
begin
  

end


endmodule