// fully-connected layer

module fc(
    input clk,

    input 
)

endmodule
