`timescale 1ns / 1ps
// memory size 30*30

module mem30x30#(parameter WIDTH = 9)
(
    input clk,
    input rst_n,
    input enable,

    input [WIDTH-1:0] data_in,

    output [WIDTH-1:0] data_out
);

// memory
reg [WIDTH-1:0] a00 [29:0];
reg [WIDTH-1:0] a01 [29:0];
reg [WIDTH-1:0] a02 [29:0];
reg [WIDTH-1:0] a03 [29:0];
reg [WIDTH-1:0] a04 [29:0];
reg [WIDTH-1:0] a05 [29:0];
reg [WIDTH-1:0] a06 [29:0];
reg [WIDTH-1:0] a07 [29:0];
reg [WIDTH-1:0] a08 [29:0];
reg [WIDTH-1:0] a09 [29:0];
reg [WIDTH-1:0] a10 [29:0];
reg [WIDTH-1:0] a11 [29:0];
reg [WIDTH-1:0] a12 [29:0];
reg [WIDTH-1:0] a13 [29:0];
reg [WIDTH-1:0] a14 [29:0];
reg [WIDTH-1:0] a15 [29:0];
reg [WIDTH-1:0] a16 [29:0];
reg [WIDTH-1:0] a17 [29:0];
reg [WIDTH-1:0] a18 [29:0];
reg [WIDTH-1:0] a19 [29:0];
reg [WIDTH-1:0] a20 [29:0];
reg [WIDTH-1:0] a21 [29:0];
reg [WIDTH-1:0] a22 [29:0];
reg [WIDTH-1:0] a23 [29:0];
reg [WIDTH-1:0] a24 [29:0];
reg [WIDTH-1:0] a25 [29:0];
reg [WIDTH-1:0] a26 [29:0];
reg [WIDTH-1:0] a27 [29:0];
reg [WIDTH-1:0] a28 [29:0];
reg [WIDTH-1:0] a29 [29:0];
// clock counter
reg [9:0] clk_counter;

// initial
initial
begin
    a00[0] <= 0;a00[1] <= 0;a00[2] <= 0;a00[3] <= 0;a00[4] <= 0;a00[5] <= 0;a00[6] <= 0;a00[7] <= 0;a00[8] <= 0;a00[9] <= 0;
    a00[10] <= 0;a00[11] <= 0;a00[12] <= 0;a00[13] <= 0;a00[14] <= 0;a00[15] <= 0;a00[16] <= 0;a00[17] <= 0;a00[18] <= 0;a00[19] <= 0;
    a00[20] <= 0;a00[21] <= 0;a00[22] <= 0;a00[23] <= 0;a00[24] <= 0;a00[25] <= 0;a00[26] <= 0;a00[27] <= 0;a00[28] <= 0;a00[29] <= 0;

    a01[0] <= 0;a01[1] <= 0;a01[2] <= 0;a01[3] <= 0;a01[4] <= 0;a01[5] <= 0;a01[6] <= 0;a01[7] <= 0;a01[8] <= 0;a01[9] <= 0;
    a01[10] <= 0;a01[11] <= 0;a01[12] <= 0;a01[13] <= 0;a01[14] <= 0;a01[15] <= 0;a01[16] <= 0;a01[17] <= 0;a01[18] <= 0;a01[19] <= 0;
    a01[20] <= 0;a01[21] <= 0;a01[22] <= 0;a01[23] <= 0;a01[24] <= 0;a01[25] <= 0;a01[26] <= 0;a01[27] <= 0;a01[28] <= 0;a01[29] <= 0;

    a02[0] <= 0;a02[1] <= 0;a02[2] <= 0;a02[3] <= 0;a02[4] <= 0;a02[5] <= 0;a02[6] <= 0;a02[7] <= 0;a02[8] <= 0;a02[9] <= 0;
    a02[10] <= 0;a02[11] <= 0;a02[12] <= 0;a02[13] <= 0;a02[14] <= 0;a02[15] <= 0;a02[16] <= 0;a02[17] <= 0;a02[18] <= 0;a02[19] <= 0;
    a02[20] <= 0;a02[21] <= 0;a02[22] <= 0;a02[23] <= 0;a02[24] <= 0;a02[25] <= 0;a02[26] <= 0;a02[27] <= 0;a02[28] <= 0;a02[29] <= 0;

	a03[0] <= 0;a03[1] <= 0;a03[2] <= 0;a03[3] <= 0;a03[4] <= 0;a03[5] <= 0;a03[6] <= 0;a03[7] <= 0;a03[8] <= 0;a03[9] <= 0;
    a03[10] <= 0;a03[11] <= 0;a03[12] <= 0;a03[13] <= 0;a03[14] <= 0;a03[15] <= 0;a03[16] <= 0;a03[17] <= 0;a03[18] <= 0;a03[19] <= 0;
    a03[20] <= 0;a03[21] <= 0;a03[22] <= 0;a03[23] <= 0;a03[24] <= 0;a03[25] <= 0;a03[26] <= 0;a03[27] <= 0;a03[28] <= 0;a03[29] <= 0;

	a04[0] <= 0;a04[1] <= 0;a04[2] <= 0;a04[3] <= 0;a04[4] <= 0;a04[5] <= 0;a04[6] <= 0;a04[7] <= 0;a04[8] <= 0;a04[9] <= 0;
    a04[10] <= 0;a04[11] <= 0;a04[12] <= 0;a04[13] <= 0;a04[14] <= 0;a04[15] <= 0;a04[16] <= 0;a04[17] <= 0;a04[18] <= 0;a04[19] <= 0;
    a04[20] <= 0;a04[21] <= 0;a04[22] <= 0;a04[23] <= 0;a04[24] <= 0;a04[25] <= 0;a04[26] <= 0;a04[27] <= 0;a04[28] <= 0;a04[29] <= 0;

	a05[0] <= 0;a05[1] <= 0;a05[2] <= 0;a05[3] <= 0;a05[4] <= 0;a05[5] <= 0;a05[6] <= 0;a05[7] <= 0;a05[8] <= 0;a05[9] <= 0;
    a05[10] <= 0;a05[11] <= 0;a05[12] <= 0;a05[13] <= 0;a05[14] <= 0;a05[15] <= 0;a05[16] <= 0;a05[17] <= 0;a05[18] <= 0;a05[19] <= 0;
    a05[20] <= 0;a05[21] <= 0;a05[22] <= 0;a05[23] <= 0;a05[24] <= 0;a05[25] <= 0;a05[26] <= 0;a05[27] <= 0;a05[28] <= 0;a05[29] <= 0;

	a06[0] <= 0;a06[1] <= 0;a06[2] <= 0;a06[3] <= 0;a06[4] <= 0;a06[5] <= 0;a06[6] <= 0;a06[7] <= 0;a06[8] <= 0;a06[9] <= 0;
    a06[10] <= 0;a06[11] <= 0;a06[12] <= 0;a06[13] <= 0;a06[14] <= 0;a06[15] <= 0;a06[16] <= 0;a06[17] <= 0;a06[18] <= 0;a06[19] <= 0;
    a06[20] <= 0;a06[21] <= 0;a06[22] <= 0;a06[23] <= 0;a06[24] <= 0;a06[25] <= 0;a06[26] <= 0;a06[27] <= 0;a06[28] <= 0;a06[29] <= 0;

    a07[0] <= 0;a07[1] <= 0;a07[2] <= 0;a07[3] <= 0;a07[4] <= 0;a07[5] <= 0;a07[6] <= 0;a07[7] <= 0;a07[8] <= 0;a07[9] <= 0;
    a07[10] <= 0;a07[11] <= 0;a07[12] <= 0;a07[13] <= 0;a07[14] <= 0;a07[15] <= 0;a07[16] <= 0;a07[17] <= 0;a07[18] <= 0;a07[19] <= 0;
    a07[20] <= 0;a07[21] <= 0;a07[22] <= 0;a07[23] <= 0;a07[24] <= 0;a07[25] <= 0;a07[26] <= 0;a07[27] <= 0;a07[28] <= 0;a07[29] <= 0;

    a08[0] <= 0;a08[1] <= 0;a08[2] <= 0;a08[3] <= 0;a08[4] <= 0;a08[5] <= 0;a08[6] <= 0;a08[7] <= 0;a08[8] <= 0;a08[9] <= 0;
    a08[10] <= 0;a08[11] <= 0;a08[12] <= 0;a08[13] <= 0;a08[14] <= 0;a08[15] <= 0;a08[16] <= 0;a08[17] <= 0;a08[18] <= 0;a08[19] <= 0;
    a08[20] <= 0;a08[21] <= 0;a08[22] <= 0;a08[23] <= 0;a08[24] <= 0;a08[25] <= 0;a08[26] <= 0;a08[27] <= 0;a08[28] <= 0;a08[29] <= 0;

    a09[0] <= 0;a09[1] <= 0;a09[2] <= 0;a09[3] <= 0;a09[4] <= 0;a09[5] <= 0;a09[6] <= 0;a09[7] <= 0;a09[8] <= 0;a09[9] <= 0;
    a09[10] <= 0;a09[11] <= 0;a09[12] <= 0;a09[13] <= 0;a09[14] <= 0;a09[15] <= 0;a09[16] <= 0;a09[17] <= 0;a09[18] <= 0;a09[19] <= 0;
    a09[20] <= 0;a09[21] <= 0;a09[22] <= 0;a09[23] <= 0;a09[24] <= 0;a09[25] <= 0;a09[26] <= 0;a09[27] <= 0;a09[28] <= 0;a09[29] <= 0;

    a10[0] <= 0;a10[1] <= 0;a10[2] <= 0;a10[3] <= 0;a10[4] <= 0;a10[5] <= 0;a10[6] <= 0;a10[7] <= 0;a10[8] <= 0;a10[9] <= 0;
    a10[10] <= 0;a10[11] <= 0;a10[12] <= 0;a10[13] <= 0;a10[14] <= 0;a10[15] <= 0;a10[16] <= 0;a10[17] <= 0;a10[18] <= 0;a10[19] <= 0;
    a10[20] <= 0;a10[21] <= 0;a10[22] <= 0;a10[23] <= 0;a10[24] <= 0;a10[25] <= 0;a10[26] <= 0;a10[27] <= 0;a10[28] <= 0;a10[29] <= 0;

    a11[0] <= 0;a11[1] <= 0;a11[2] <= 0;a11[3] <= 0;a11[4] <= 0;a11[5] <= 0;a11[6] <= 0;a11[7] <= 0;a11[8] <= 0;a11[9] <= 0;
    a11[10] <= 0;a11[11] <= 0;a11[12] <= 0;a11[13] <= 0;a11[14] <= 0;a11[15] <= 0;a11[16] <= 0;a11[17] <= 0;a11[18] <= 0;a11[19] <= 0;
    a11[20] <= 0;a11[21] <= 0;a11[22] <= 0;a11[23] <= 0;a11[24] <= 0;a11[25] <= 0;a11[26] <= 0;a11[27] <= 0;a11[28] <= 0;a11[29] <= 0;

    a12[0] <= 0;a12[1] <= 0;a12[2] <= 0;a12[3] <= 0;a12[4] <= 0;a12[5] <= 0;a12[6] <= 0;a12[7] <= 0;a12[8] <= 0;a12[9] <= 0;
    a12[10] <= 0;a12[11] <= 0;a12[12] <= 0;a12[13] <= 0;a12[14] <= 0;a12[15] <= 0;a12[16] <= 0;a12[17] <= 0;a12[18] <= 0;a12[19] <= 0;
    a12[20] <= 0;a12[21] <= 0;a12[22] <= 0;a12[23] <= 0;a12[24] <= 0;a12[25] <= 0;a12[26] <= 0;a12[27] <= 0;a12[28] <= 0;a12[29] <= 0;

    a13[0] <= 0;a13[1] <= 0;a13[2] <= 0;a13[3] <= 0;a13[4] <= 0;a13[5] <= 0;a13[6] <= 0;a13[7] <= 0;a13[8] <= 0;a13[9] <= 0;
    a13[10] <= 0;a13[11] <= 0;a13[12] <= 0;a13[13] <= 0;a13[14] <= 0;a13[15] <= 0;a13[16] <= 0;a13[17] <= 0;a13[18] <= 0;a13[19] <= 0;
    a13[20] <= 0;a13[21] <= 0;a13[22] <= 0;a13[23] <= 0;a13[24] <= 0;a13[25] <= 0;a13[26] <= 0;a13[27] <= 0;a13[28] <= 0;a13[29] <= 0;

    a14[0] <= 0;a14[1] <= 0;a14[2] <= 0;a14[3] <= 0;a14[4] <= 0;a14[5] <= 0;a14[6] <= 0;a14[7] <= 0;a14[8] <= 0;a14[9] <= 0;
    a14[10] <= 0;a14[11] <= 0;a14[12] <= 0;a14[13] <= 0;a14[14] <= 0;a14[15] <= 0;a14[16] <= 0;a14[17] <= 0;a14[18] <= 0;a14[19] <= 0;
    a14[20] <= 0;a14[21] <= 0;a14[22] <= 0;a14[23] <= 0;a14[24] <= 0;a14[25] <= 0;a14[26] <= 0;a14[27] <= 0;a14[28] <= 0;a14[29] <= 0;

    a15[0] <= 0;a15[1] <= 0;a15[2] <= 0;a15[3] <= 0;a15[4] <= 0;a15[5] <= 0;a15[6] <= 0;a15[7] <= 0;a15[8] <= 0;a15[9] <= 0;
    a15[10] <= 0;a15[11] <= 0;a15[12] <= 0;a15[13] <= 0;a15[14] <= 0;a15[15] <= 0;a15[16] <= 0;a15[17] <= 0;a15[18] <= 0;a15[19] <= 0;
    a15[20] <= 0;a15[21] <= 0;a15[22] <= 0;a15[23] <= 0;a15[24] <= 0;a15[25] <= 0;a15[26] <= 0;a15[27] <= 0;a15[28] <= 0;a15[29] <= 0;

    a16[0] <= 0;a16[1] <= 0;a16[2] <= 0;a16[3] <= 0;a16[4] <= 0;a16[5] <= 0;a16[6] <= 0;a16[7] <= 0;a16[8] <= 0;a16[9] <= 0;
    a16[10] <= 0;a16[11] <= 0;a16[12] <= 0;a16[13] <= 0;a16[14] <= 0;a16[15] <= 0;a16[16] <= 0;a16[17] <= 0;a16[18] <= 0;a16[19] <= 0;
    a16[20] <= 0;a16[21] <= 0;a16[22] <= 0;a16[23] <= 0;a16[24] <= 0;a16[25] <= 0;a16[26] <= 0;a16[27] <= 0;a16[28] <= 0;a16[29] <= 0;

    a17[0] <= 0;a17[1] <= 0;a17[2] <= 0;a17[3] <= 0;a17[4] <= 0;a17[5] <= 0;a17[6] <= 0;a17[7] <= 0;a17[8] <= 0;a17[9] <= 0;
    a17[10] <= 0;a17[11] <= 0;a17[12] <= 0;a17[13] <= 0;a17[14] <= 0;a17[15] <= 0;a17[16] <= 0;a17[17] <= 0;a17[18] <= 0;a17[19] <= 0;
    a17[20] <= 0;a17[21] <= 0;a17[22] <= 0;a17[23] <= 0;a17[24] <= 0;a17[25] <= 0;a17[26] <= 0;a17[27] <= 0;a17[28] <= 0;a17[29] <= 0;

    a18[0] <= 0;a18[1] <= 0;a18[2] <= 0;a18[3] <= 0;a18[4] <= 0;a18[5] <= 0;a18[6] <= 0;a18[7] <= 0;a18[8] <= 0;a18[9] <= 0;
    a18[10] <= 0;a18[11] <= 0;a18[12] <= 0;a18[13] <= 0;a18[14] <= 0;a18[15] <= 0;a18[16] <= 0;a18[17] <= 0;a18[18] <= 0;a18[19] <= 0;
    a18[20] <= 0;a18[21] <= 0;a18[22] <= 0;a18[23] <= 0;a18[24] <= 0;a18[25] <= 0;a18[26] <= 0;a18[27] <= 0;a18[28] <= 0;a18[29] <= 0;

    a19[0] <= 0;a19[1] <= 0;a19[2] <= 0;a19[3] <= 0;a19[4] <= 0;a19[5] <= 0;a19[6] <= 0;a19[7] <= 0;a19[8] <= 0;a19[9] <= 0;
    a19[10] <= 0;a19[11] <= 0;a19[12] <= 0;a19[13] <= 0;a19[14] <= 0;a19[15] <= 0;a19[16] <= 0;a19[17] <= 0;a19[18] <= 0;a19[19] <= 0;
    a19[20] <= 0;a19[21] <= 0;a19[22] <= 0;a19[23] <= 0;a19[24] <= 0;a19[25] <= 0;a19[26] <= 0;a19[27] <= 0;a19[28] <= 0;a19[29] <= 0;

    a20[0] <= 0;a20[1] <= 0;a20[2] <= 0;a20[3] <= 0;a20[4] <= 0;a20[5] <= 0;a20[6] <= 0;a20[7] <= 0;a20[8] <= 0;a20[9] <= 0;
    a20[10] <= 0;a20[11] <= 0;a20[12] <= 0;a20[13] <= 0;a20[14] <= 0;a20[15] <= 0;a20[16] <= 0;a20[17] <= 0;a20[18] <= 0;a20[19] <= 0;
    a20[20] <= 0;a20[21] <= 0;a20[22] <= 0;a20[23] <= 0;a20[24] <= 0;a20[25] <= 0;a20[26] <= 0;a20[27] <= 0;a20[28] <= 0;a20[29] <= 0;

    a21[0] <= 0;a21[1] <= 0;a21[2] <= 0;a21[3] <= 0;a21[4] <= 0;a21[5] <= 0;a21[6] <= 0;a21[7] <= 0;a21[8] <= 0;a21[9] <= 0;
    a21[10] <= 0;a21[11] <= 0;a21[12] <= 0;a21[13] <= 0;a21[14] <= 0;a21[15] <= 0;a21[16] <= 0;a21[17] <= 0;a21[18] <= 0;a21[19] <= 0;
    a21[20] <= 0;a21[21] <= 0;a21[22] <= 0;a21[23] <= 0;a21[24] <= 0;a21[25] <= 0;a21[26] <= 0;a21[27] <= 0;a21[28] <= 0;a21[29] <= 0;

    a22[0] <= 0;a22[1] <= 0;a22[2] <= 0;a22[3] <= 0;a22[4] <= 0;a22[5] <= 0;a22[6] <= 0;a22[7] <= 0;a22[8] <= 0;a22[9] <= 0;
    a22[10] <= 0;a22[11] <= 0;a22[12] <= 0;a22[13] <= 0;a22[14] <= 0;a22[15] <= 0;a22[16] <= 0;a22[17] <= 0;a22[18] <= 0;a22[19] <= 0;
    a22[20] <= 0;a22[21] <= 0;a22[22] <= 0;a22[23] <= 0;a22[24] <= 0;a22[25] <= 0;a22[26] <= 0;a22[27] <= 0;a22[28] <= 0;a22[29] <= 0;

    a23[0] <= 0;a23[1] <= 0;a23[2] <= 0;a23[3] <= 0;a23[4] <= 0;a23[5] <= 0;a23[6] <= 0;a23[7] <= 0;a23[8] <= 0;a23[9] <= 0;
    a23[10] <= 0;a23[11] <= 0;a23[12] <= 0;a23[13] <= 0;a23[14] <= 0;a23[15] <= 0;a23[16] <= 0;a23[17] <= 0;a23[18] <= 0;a23[19] <= 0;
    a23[20] <= 0;a23[21] <= 0;a23[22] <= 0;a23[23] <= 0;a23[24] <= 0;a23[25] <= 0;a23[26] <= 0;a23[27] <= 0;a23[28] <= 0;a23[29] <= 0;

    a24[0] <= 0;a24[1] <= 0;a24[2] <= 0;a24[3] <= 0;a24[4] <= 0;a24[5] <= 0;a24[6] <= 0;a24[7] <= 0;a24[8] <= 0;a24[9] <= 0;
    a24[10] <= 0;a24[11] <= 0;a24[12] <= 0;a24[13] <= 0;a24[14] <= 0;a24[15] <= 0;a24[16] <= 0;a24[17] <= 0;a24[18] <= 0;a24[19] <= 0;
    a24[20] <= 0;a24[21] <= 0;a24[22] <= 0;a24[23] <= 0;a24[24] <= 0;a24[25] <= 0;a24[26] <= 0;a24[27] <= 0;a24[28] <= 0;a24[29] <= 0;

    a25[0] <= 0;a25[1] <= 0;a25[2] <= 0;a25[3] <= 0;a25[4] <= 0;a25[5] <= 0;a25[6] <= 0;a25[7] <= 0;a25[8] <= 0;a25[9] <= 0;
    a25[10] <= 0;a25[11] <= 0;a25[12] <= 0;a25[13] <= 0;a25[14] <= 0;a25[15] <= 0;a25[16] <= 0;a25[17] <= 0;a25[18] <= 0;a25[19] <= 0;
    a25[20] <= 0;a25[21] <= 0;a25[22] <= 0;a25[23] <= 0;a25[24] <= 0;a25[25] <= 0;a25[26] <= 0;a25[27] <= 0;a25[28] <= 0;a25[29] <= 0;

    a26[0] <= 0;a26[1] <= 0;a26[2] <= 0;a26[3] <= 0;a26[4] <= 0;a26[5] <= 0;a26[6] <= 0;a26[7] <= 0;a26[8] <= 0;a26[9] <= 0;
    a26[10] <= 0;a26[11] <= 0;a26[12] <= 0;a26[13] <= 0;a26[14] <= 0;a26[15] <= 0;a26[16] <= 0;a26[17] <= 0;a26[18] <= 0;a26[19] <= 0;
    a26[20] <= 0;a26[21] <= 0;a26[22] <= 0;a26[23] <= 0;a26[24] <= 0;a26[25] <= 0;a26[26] <= 0;a26[27] <= 0;a26[28] <= 0;a26[29] <= 0;

    a27[0] <= 0;a27[1] <= 0;a27[2] <= 0;a27[3] <= 0;a27[4] <= 0;a27[5] <= 0;a27[6] <= 0;a27[7] <= 0;a27[8] <= 0;a27[9] <= 0;
    a27[10] <= 0;a27[11] <= 0;a27[12] <= 0;a27[13] <= 0;a27[14] <= 0;a27[15] <= 0;a27[16] <= 0;a27[17] <= 0;a27[18] <= 0;a27[19] <= 0;
    a27[20] <= 0;a27[21] <= 0;a27[22] <= 0;a27[23] <= 0;a27[24] <= 0;a27[25] <= 0;a27[26] <= 0;a27[27] <= 0;a27[28] <= 0;a27[29] <= 0;

    a28[0] <= 0;a28[1] <= 0;a28[2] <= 0;a28[3] <= 0;a28[4] <= 0;a28[5] <= 0;a28[6] <= 0;a28[7] <= 0;a28[8] <= 0;a28[9] <= 0;
    a28[10] <= 0;a28[11] <= 0;a28[12] <= 0;a28[13] <= 0;a28[14] <= 0;a28[15] <= 0;a28[16] <= 0;a28[17] <= 0;a28[18] <= 0;a28[19] <= 0;
    a28[20] <= 0;a28[21] <= 0;a28[22] <= 0;a28[23] <= 0;a28[24] <= 0;a28[25] <= 0;a28[26] <= 0;a28[27] <= 0;a28[28] <= 0;a28[29] <= 0;

    a29[0] <= 0;a29[1] <= 0;a29[2] <= 0;a29[3] <= 0;a29[4] <= 0;a29[5] <= 0;a29[6] <= 0;a29[7] <= 0;a29[8] <= 0;a29[9] <= 0;
    a29[10] <= 0;a29[11] <= 0;a29[12] <= 0;a29[13] <= 0;a29[14] <= 0;a29[15] <= 0;a29[16] <= 0;a29[17] <= 0;a29[18] <= 0;a29[19] <= 0;
    a29[20] <= 0;a29[21] <= 0;a29[22] <= 0;a29[23] <= 0;a29[24] <= 0;a29[25] <= 0;a29[26] <= 0;a29[27] <= 0;a29[28] <= 0;a29[29] <= 0;

    clk_counter = 0;
end

always@(posedge clk)
begin
    if((!rst_n)&&enable)
    begin
        a00[0] <= data_in;
        case (clk_counter)
            0:
			begin
				a00[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			1:
			begin
				a00[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			2:
			begin
				a00[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			3:
			begin
				a00[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			4:
			begin
				a00[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			5:
			begin
				a00[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			6:
			begin
				a00[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			7:
			begin
				a00[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			8:
			begin
				a00[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			9:
			begin
				a00[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			10:
			begin
				a00[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			11:
			begin
				a00[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			12:
			begin
				a00[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			13:
			begin
				a00[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			14:
			begin
				a00[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			15:
			begin
				a00[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			16:
			begin
				a00[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			17:
			begin
				a00[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			18:
			begin
				a00[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			19:
			begin
				a00[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			20:
			begin
				a00[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			21:
			begin
				a00[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			22:
			begin
				a00[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			23:
			begin
				a00[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			24:
			begin
				a00[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			25:
			begin
				a00[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			26:
			begin
				a00[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			27:
			begin
				a00[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			28:
			begin
				a00[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			29:
			begin
				a00[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			30:
			begin
				a01[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			31:
			begin
				a01[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			32:
			begin
				a01[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			33:
			begin
				a01[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			34:
			begin
				a01[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			35:
			begin
				a01[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			36:
			begin
				a01[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			37:
			begin
				a01[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			38:
			begin
				a01[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			39:
			begin
				a01[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			40:
			begin
				a01[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			41:
			begin
				a01[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			42:
			begin
				a01[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			43:
			begin
				a01[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			44:
			begin
				a01[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			45:
			begin
				a01[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			46:
			begin
				a01[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			47:
			begin
				a01[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			48:
			begin
				a01[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			49:
			begin
				a01[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			50:
			begin
				a01[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			51:
			begin
				a01[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			52:
			begin
				a01[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			53:
			begin
				a01[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			54:
			begin
				a01[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			55:
			begin
				a01[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			56:
			begin
				a01[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			57:
			begin
				a01[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			58:
			begin
				a01[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			59:
			begin
				a01[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			60:
			begin
				a02[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			61:
			begin
				a02[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			62:
			begin
				a02[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			63:
			begin
				a02[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			64:
			begin
				a02[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			65:
			begin
				a02[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			66:
			begin
				a02[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			67:
			begin
				a02[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			68:
			begin
				a02[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			69:
			begin
				a02[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			70:
			begin
				a02[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			71:
			begin
				a02[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			72:
			begin
				a02[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			73:
			begin
				a02[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			74:
			begin
				a02[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			75:
			begin
				a02[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			76:
			begin
				a02[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			77:
			begin
				a02[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			78:
			begin
				a02[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			79:
			begin
				a02[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			80:
			begin
				a02[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			81:
			begin
				a02[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			82:
			begin
				a02[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			83:
			begin
				a02[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			84:
			begin
				a02[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			85:
			begin
				a02[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			86:
			begin
				a02[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			87:
			begin
				a02[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			88:
			begin
				a02[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			89:
			begin
				a02[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			90:
			begin
				a03[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			91:
			begin
				a03[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			92:
			begin
				a03[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			93:
			begin
				a03[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			94:
			begin
				a03[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			95:
			begin
				a03[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			96:
			begin
				a03[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			97:
			begin
				a03[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			98:
			begin
				a03[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			99:
			begin
				a03[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			100:
			begin
				a03[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			101:
			begin
				a03[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			102:
			begin
				a03[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			103:
			begin
				a03[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			104:
			begin
				a03[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			105:
			begin
				a03[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			106:
			begin
				a03[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			107:
			begin
				a03[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			108:
			begin
				a03[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			109:
			begin
				a03[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			110:
			begin
				a03[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			111:
			begin
				a03[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			112:
			begin
				a03[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			113:
			begin
				a03[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			114:
			begin
				a03[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			115:
			begin
				a03[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			116:
			begin
				a03[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			117:
			begin
				a03[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			118:
			begin
				a03[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			119:
			begin
				a03[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			120:
			begin
				a04[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			121:
			begin
				a04[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			122:
			begin
				a04[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			123:
			begin
				a04[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			124:
			begin
				a04[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			125:
			begin
				a04[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			126:
			begin
				a04[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			127:
			begin
				a04[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			128:
			begin
				a04[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			129:
			begin
				a04[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			130:
			begin
				a04[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			131:
			begin
				a04[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			132:
			begin
				a04[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			133:
			begin
				a04[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			134:
			begin
				a04[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			135:
			begin
				a04[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			136:
			begin
				a04[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			137:
			begin
				a04[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			138:
			begin
				a04[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			139:
			begin
				a04[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			140:
			begin
				a04[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			141:
			begin
				a04[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			142:
			begin
				a04[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			143:
			begin
				a04[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			144:
			begin
				a04[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			145:
			begin
				a04[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			146:
			begin
				a04[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			147:
			begin
				a04[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			148:
			begin
				a04[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			149:
			begin
				a04[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			150:
			begin
				a05[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			151:
			begin
				a05[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			152:
			begin
				a05[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			153:
			begin
				a05[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			154:
			begin
				a05[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			155:
			begin
				a05[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			156:
			begin
				a05[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			157:
			begin
				a05[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			158:
			begin
				a05[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			159:
			begin
				a05[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			160:
			begin
				a05[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			161:
			begin
				a05[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			162:
			begin
				a05[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			163:
			begin
				a05[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			164:
			begin
				a05[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			165:
			begin
				a05[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			166:
			begin
				a05[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			167:
			begin
				a05[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			168:
			begin
				a05[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			169:
			begin
				a05[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			170:
			begin
				a05[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			171:
			begin
				a05[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			172:
			begin
				a05[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			173:
			begin
				a05[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			174:
			begin
				a05[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			175:
			begin
				a05[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			176:
			begin
				a05[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			177:
			begin
				a05[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			178:
			begin
				a05[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			179:
			begin
				a05[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			180:
			begin
				a06[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			181:
			begin
				a06[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			182:
			begin
				a06[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			183:
			begin
				a06[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			184:
			begin
				a06[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			185:
			begin
				a06[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			186:
			begin
				a06[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			187:
			begin
				a06[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			188:
			begin
				a06[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			189:
			begin
				a06[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			190:
			begin
				a06[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			191:
			begin
				a06[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			192:
			begin
				a06[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			193:
			begin
				a06[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			194:
			begin
				a06[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			195:
			begin
				a06[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			196:
			begin
				a06[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			197:
			begin
				a06[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			198:
			begin
				a06[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			199:
			begin
				a06[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			200:
			begin
				a06[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			201:
			begin
				a06[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			202:
			begin
				a06[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			203:
			begin
				a06[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			204:
			begin
				a06[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			205:
			begin
				a06[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			206:
			begin
				a06[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			207:
			begin
				a06[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			208:
			begin
				a06[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			209:
			begin
				a06[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			210:
			begin
				a07[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			211:
			begin
				a07[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			212:
			begin
				a07[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			213:
			begin
				a07[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			214:
			begin
				a07[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			215:
			begin
				a07[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			216:
			begin
				a07[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			217:
			begin
				a07[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			218:
			begin
				a07[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			219:
			begin
				a07[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			220:
			begin
				a07[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			221:
			begin
				a07[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			222:
			begin
				a07[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			223:
			begin
				a07[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			224:
			begin
				a07[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			225:
			begin
				a07[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			226:
			begin
				a07[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			227:
			begin
				a07[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			228:
			begin
				a07[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			229:
			begin
				a07[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			230:
			begin
				a07[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			231:
			begin
				a07[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			232:
			begin
				a07[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			233:
			begin
				a07[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			234:
			begin
				a07[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			235:
			begin
				a07[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			236:
			begin
				a07[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			237:
			begin
				a07[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			238:
			begin
				a07[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			239:
			begin
				a07[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			240:
			begin
				a08[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			241:
			begin
				a08[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			242:
			begin
				a08[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			243:
			begin
				a08[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			244:
			begin
				a08[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			245:
			begin
				a08[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			246:
			begin
				a08[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			247:
			begin
				a08[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			248:
			begin
				a08[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			249:
			begin
				a08[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			250:
			begin
				a08[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			251:
			begin
				a08[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			252:
			begin
				a08[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			253:
			begin
				a08[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			254:
			begin
				a08[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			255:
			begin
				a08[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			256:
			begin
				a08[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			257:
			begin
				a08[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			258:
			begin
				a08[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			259:
			begin
				a08[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			260:
			begin
				a08[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			261:
			begin
				a08[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			262:
			begin
				a08[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			263:
			begin
				a08[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			264:
			begin
				a08[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			265:
			begin
				a08[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			266:
			begin
				a08[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			267:
			begin
				a08[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			268:
			begin
				a08[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			269:
			begin
				a08[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			270:
			begin
				a09[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			271:
			begin
				a09[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			272:
			begin
				a09[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			273:
			begin
				a09[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			274:
			begin
				a09[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			275:
			begin
				a09[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			276:
			begin
				a09[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			277:
			begin
				a09[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			278:
			begin
				a09[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			279:
			begin
				a09[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			280:
			begin
				a09[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			281:
			begin
				a09[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			282:
			begin
				a09[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			283:
			begin
				a09[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			284:
			begin
				a09[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			285:
			begin
				a09[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			286:
			begin
				a09[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			287:
			begin
				a09[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			288:
			begin
				a09[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			289:
			begin
				a09[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			290:
			begin
				a09[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			291:
			begin
				a09[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			292:
			begin
				a09[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			293:
			begin
				a09[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			294:
			begin
				a09[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			295:
			begin
				a09[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			296:
			begin
				a09[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			297:
			begin
				a09[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			298:
			begin
				a09[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			299:
			begin
				a09[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			300:
			begin
				a10[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			301:
			begin
				a10[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			302:
			begin
				a10[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			303:
			begin
				a10[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			304:
			begin
				a10[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			305:
			begin
				a10[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			306:
			begin
				a10[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			307:
			begin
				a10[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			308:
			begin
				a10[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			309:
			begin
				a10[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			310:
			begin
				a10[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			311:
			begin
				a10[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			312:
			begin
				a10[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			313:
			begin
				a10[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			314:
			begin
				a10[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			315:
			begin
				a10[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			316:
			begin
				a10[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			317:
			begin
				a10[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			318:
			begin
				a10[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			319:
			begin
				a10[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			320:
			begin
				a10[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			321:
			begin
				a10[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			322:
			begin
				a10[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			323:
			begin
				a10[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			324:
			begin
				a10[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			325:
			begin
				a10[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			326:
			begin
				a10[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			327:
			begin
				a10[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			328:
			begin
				a10[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			329:
			begin
				a10[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			330:
			begin
				a11[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			331:
			begin
				a11[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			332:
			begin
				a11[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			333:
			begin
				a11[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			334:
			begin
				a11[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			335:
			begin
				a11[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			336:
			begin
				a11[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			337:
			begin
				a11[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			338:
			begin
				a11[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			339:
			begin
				a11[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			340:
			begin
				a11[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			341:
			begin
				a11[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			342:
			begin
				a11[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			343:
			begin
				a11[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			344:
			begin
				a11[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			345:
			begin
				a11[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			346:
			begin
				a11[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			347:
			begin
				a11[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			348:
			begin
				a11[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			349:
			begin
				a11[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			350:
			begin
				a11[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			351:
			begin
				a11[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			352:
			begin
				a11[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			353:
			begin
				a11[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			354:
			begin
				a11[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			355:
			begin
				a11[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			356:
			begin
				a11[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			357:
			begin
				a11[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			358:
			begin
				a11[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			359:
			begin
				a11[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			360:
			begin
				a12[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			361:
			begin
				a12[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			362:
			begin
				a12[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			363:
			begin
				a12[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			364:
			begin
				a12[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			365:
			begin
				a12[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			366:
			begin
				a12[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			367:
			begin
				a12[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			368:
			begin
				a12[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			369:
			begin
				a12[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			370:
			begin
				a12[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			371:
			begin
				a12[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			372:
			begin
				a12[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			373:
			begin
				a12[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			374:
			begin
				a12[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			375:
			begin
				a12[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			376:
			begin
				a12[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			377:
			begin
				a12[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			378:
			begin
				a12[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			379:
			begin
				a12[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			380:
			begin
				a12[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			381:
			begin
				a12[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			382:
			begin
				a12[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			383:
			begin
				a12[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			384:
			begin
				a12[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			385:
			begin
				a12[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			386:
			begin
				a12[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			387:
			begin
				a12[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			388:
			begin
				a12[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			389:
			begin
				a12[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			390:
			begin
				a13[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			391:
			begin
				a13[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			392:
			begin
				a13[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			393:
			begin
				a13[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			394:
			begin
				a13[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			395:
			begin
				a13[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			396:
			begin
				a13[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			397:
			begin
				a13[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			398:
			begin
				a13[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			399:
			begin
				a13[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			400:
			begin
				a13[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			401:
			begin
				a13[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			402:
			begin
				a13[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			403:
			begin
				a13[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			404:
			begin
				a13[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			405:
			begin
				a13[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			406:
			begin
				a13[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			407:
			begin
				a13[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			408:
			begin
				a13[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			409:
			begin
				a13[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			410:
			begin
				a13[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			411:
			begin
				a13[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			412:
			begin
				a13[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			413:
			begin
				a13[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			414:
			begin
				a13[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			415:
			begin
				a13[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			416:
			begin
				a13[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			417:
			begin
				a13[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			418:
			begin
				a13[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			419:
			begin
				a13[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			420:
			begin
				a14[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			421:
			begin
				a14[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			422:
			begin
				a14[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			423:
			begin
				a14[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			424:
			begin
				a14[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			425:
			begin
				a14[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			426:
			begin
				a14[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			427:
			begin
				a14[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			428:
			begin
				a14[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			429:
			begin
				a14[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			430:
			begin
				a14[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			431:
			begin
				a14[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			432:
			begin
				a14[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			433:
			begin
				a14[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			434:
			begin
				a14[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			435:
			begin
				a14[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			436:
			begin
				a14[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			437:
			begin
				a14[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			438:
			begin
				a14[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			439:
			begin
				a14[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			440:
			begin
				a14[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			441:
			begin
				a14[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			442:
			begin
				a14[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			443:
			begin
				a14[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			444:
			begin
				a14[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			445:
			begin
				a14[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			446:
			begin
				a14[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			447:
			begin
				a14[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			448:
			begin
				a14[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			449:
			begin
				a14[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			450:
			begin
				a15[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			451:
			begin
				a15[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			452:
			begin
				a15[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			453:
			begin
				a15[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			454:
			begin
				a15[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			455:
			begin
				a15[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			456:
			begin
				a15[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			457:
			begin
				a15[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			458:
			begin
				a15[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			459:
			begin
				a15[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			460:
			begin
				a15[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			461:
			begin
				a15[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			462:
			begin
				a15[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			463:
			begin
				a15[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			464:
			begin
				a15[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			465:
			begin
				a15[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			466:
			begin
				a15[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			467:
			begin
				a15[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			468:
			begin
				a15[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			469:
			begin
				a15[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			470:
			begin
				a15[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			471:
			begin
				a15[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			472:
			begin
				a15[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			473:
			begin
				a15[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			474:
			begin
				a15[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			475:
			begin
				a15[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			476:
			begin
				a15[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			477:
			begin
				a15[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			478:
			begin
				a15[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			479:
			begin
				a15[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			480:
			begin
				a16[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			481:
			begin
				a16[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			482:
			begin
				a16[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			483:
			begin
				a16[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			484:
			begin
				a16[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			485:
			begin
				a16[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			486:
			begin
				a16[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			487:
			begin
				a16[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			488:
			begin
				a16[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			489:
			begin
				a16[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			490:
			begin
				a16[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			491:
			begin
				a16[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			492:
			begin
				a16[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			493:
			begin
				a16[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			494:
			begin
				a16[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			495:
			begin
				a16[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			496:
			begin
				a16[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			497:
			begin
				a16[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			498:
			begin
				a16[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			499:
			begin
				a16[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			500:
			begin
				a16[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			501:
			begin
				a16[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			502:
			begin
				a16[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			503:
			begin
				a16[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			504:
			begin
				a16[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			505:
			begin
				a16[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			506:
			begin
				a16[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			507:
			begin
				a16[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			508:
			begin
				a16[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			509:
			begin
				a16[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			510:
			begin
				a17[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			511:
			begin
				a17[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			512:
			begin
				a17[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			513:
			begin
				a17[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			514:
			begin
				a17[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			515:
			begin
				a17[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			516:
			begin
				a17[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			517:
			begin
				a17[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			518:
			begin
				a17[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			519:
			begin
				a17[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			520:
			begin
				a17[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			521:
			begin
				a17[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			522:
			begin
				a17[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			523:
			begin
				a17[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			524:
			begin
				a17[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			525:
			begin
				a17[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			526:
			begin
				a17[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			527:
			begin
				a17[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			528:
			begin
				a17[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			529:
			begin
				a17[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			530:
			begin
				a17[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			531:
			begin
				a17[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			532:
			begin
				a17[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			533:
			begin
				a17[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			534:
			begin
				a17[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			535:
			begin
				a17[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			536:
			begin
				a17[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			537:
			begin
				a17[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			538:
			begin
				a17[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			539:
			begin
				a17[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			540:
			begin
				a18[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			541:
			begin
				a18[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			542:
			begin
				a18[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			543:
			begin
				a18[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			544:
			begin
				a18[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			545:
			begin
				a18[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			546:
			begin
				a18[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			547:
			begin
				a18[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			548:
			begin
				a18[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			549:
			begin
				a18[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			550:
			begin
				a18[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			551:
			begin
				a18[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			552:
			begin
				a18[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			553:
			begin
				a18[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			554:
			begin
				a18[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			555:
			begin
				a18[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			556:
			begin
				a18[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			557:
			begin
				a18[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			558:
			begin
				a18[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			559:
			begin
				a18[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			560:
			begin
				a18[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			561:
			begin
				a18[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			562:
			begin
				a18[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			563:
			begin
				a18[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			564:
			begin
				a18[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			565:
			begin
				a18[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			566:
			begin
				a18[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			567:
			begin
				a18[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			568:
			begin
				a18[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			569:
			begin
				a18[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			570:
			begin
				a19[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			571:
			begin
				a19[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			572:
			begin
				a19[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			573:
			begin
				a19[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			574:
			begin
				a19[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			575:
			begin
				a19[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			576:
			begin
				a19[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			577:
			begin
				a19[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			578:
			begin
				a19[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			579:
			begin
				a19[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			580:
			begin
				a19[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			581:
			begin
				a19[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			582:
			begin
				a19[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			583:
			begin
				a19[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			584:
			begin
				a19[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			585:
			begin
				a19[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			586:
			begin
				a19[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			587:
			begin
				a19[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			588:
			begin
				a19[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			589:
			begin
				a19[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			590:
			begin
				a19[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			591:
			begin
				a19[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			592:
			begin
				a19[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			593:
			begin
				a19[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			594:
			begin
				a19[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			595:
			begin
				a19[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			596:
			begin
				a19[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			597:
			begin
				a19[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			598:
			begin
				a19[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			599:
			begin
				a19[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			600:
			begin
				a20[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			601:
			begin
				a20[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			602:
			begin
				a20[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			603:
			begin
				a20[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			604:
			begin
				a20[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			605:
			begin
				a20[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			606:
			begin
				a20[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			607:
			begin
				a20[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			608:
			begin
				a20[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			609:
			begin
				a20[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			610:
			begin
				a20[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			611:
			begin
				a20[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			612:
			begin
				a20[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			613:
			begin
				a20[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			614:
			begin
				a20[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			615:
			begin
				a20[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			616:
			begin
				a20[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			617:
			begin
				a20[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			618:
			begin
				a20[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			619:
			begin
				a20[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			620:
			begin
				a20[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			621:
			begin
				a20[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			622:
			begin
				a20[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			623:
			begin
				a20[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			624:
			begin
				a20[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			625:
			begin
				a20[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			626:
			begin
				a20[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			627:
			begin
				a20[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			628:
			begin
				a20[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			629:
			begin
				a20[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			630:
			begin
				a21[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			631:
			begin
				a21[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			632:
			begin
				a21[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			633:
			begin
				a21[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			634:
			begin
				a21[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			635:
			begin
				a21[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			636:
			begin
				a21[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			637:
			begin
				a21[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			638:
			begin
				a21[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			639:
			begin
				a21[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			640:
			begin
				a21[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			641:
			begin
				a21[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			642:
			begin
				a21[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			643:
			begin
				a21[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			644:
			begin
				a21[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			645:
			begin
				a21[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			646:
			begin
				a21[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			647:
			begin
				a21[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			648:
			begin
				a21[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			649:
			begin
				a21[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			650:
			begin
				a21[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			651:
			begin
				a21[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			652:
			begin
				a21[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			653:
			begin
				a21[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			654:
			begin
				a21[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			655:
			begin
				a21[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			656:
			begin
				a21[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			657:
			begin
				a21[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			658:
			begin
				a21[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			659:
			begin
				a21[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			660:
			begin
				a22[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			661:
			begin
				a22[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			662:
			begin
				a22[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			663:
			begin
				a22[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			664:
			begin
				a22[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			665:
			begin
				a22[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			666:
			begin
				a22[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			667:
			begin
				a22[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			668:
			begin
				a22[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			669:
			begin
				a22[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			670:
			begin
				a22[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			671:
			begin
				a22[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			672:
			begin
				a22[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			673:
			begin
				a22[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			674:
			begin
				a22[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			675:
			begin
				a22[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			676:
			begin
				a22[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			677:
			begin
				a22[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			678:
			begin
				a22[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			679:
			begin
				a22[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			680:
			begin
				a22[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			681:
			begin
				a22[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			682:
			begin
				a22[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			683:
			begin
				a22[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			684:
			begin
				a22[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			685:
			begin
				a22[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			686:
			begin
				a22[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			687:
			begin
				a22[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			688:
			begin
				a22[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			689:
			begin
				a22[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			690:
			begin
				a23[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			691:
			begin
				a23[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			692:
			begin
				a23[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			693:
			begin
				a23[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			694:
			begin
				a23[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			695:
			begin
				a23[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			696:
			begin
				a23[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			697:
			begin
				a23[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			698:
			begin
				a23[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			699:
			begin
				a23[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			700:
			begin
				a23[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			701:
			begin
				a23[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			702:
			begin
				a23[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			703:
			begin
				a23[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			704:
			begin
				a23[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			705:
			begin
				a23[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			706:
			begin
				a23[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			707:
			begin
				a23[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			708:
			begin
				a23[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			709:
			begin
				a23[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			710:
			begin
				a23[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			711:
			begin
				a23[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			712:
			begin
				a23[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			713:
			begin
				a23[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			714:
			begin
				a23[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			715:
			begin
				a23[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			716:
			begin
				a23[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			717:
			begin
				a23[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			718:
			begin
				a23[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			719:
			begin
				a23[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			720:
			begin
				a24[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			721:
			begin
				a24[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			722:
			begin
				a24[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			723:
			begin
				a24[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			724:
			begin
				a24[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			725:
			begin
				a24[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			726:
			begin
				a24[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			727:
			begin
				a24[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			728:
			begin
				a24[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			729:
			begin
				a24[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			730:
			begin
				a24[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			731:
			begin
				a24[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			732:
			begin
				a24[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			733:
			begin
				a24[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			734:
			begin
				a24[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			735:
			begin
				a24[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			736:
			begin
				a24[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			737:
			begin
				a24[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			738:
			begin
				a24[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			739:
			begin
				a24[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			740:
			begin
				a24[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			741:
			begin
				a24[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			742:
			begin
				a24[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			743:
			begin
				a24[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			744:
			begin
				a24[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			745:
			begin
				a24[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			746:
			begin
				a24[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			747:
			begin
				a24[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			748:
			begin
				a24[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			749:
			begin
				a24[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			750:
			begin
				a25[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			751:
			begin
				a25[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			752:
			begin
				a25[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			753:
			begin
				a25[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			754:
			begin
				a25[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			755:
			begin
				a25[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			756:
			begin
				a25[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			757:
			begin
				a25[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			758:
			begin
				a25[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			759:
			begin
				a25[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			760:
			begin
				a25[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			761:
			begin
				a25[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			762:
			begin
				a25[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			763:
			begin
				a25[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			764:
			begin
				a25[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			765:
			begin
				a25[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			766:
			begin
				a25[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			767:
			begin
				a25[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			768:
			begin
				a25[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			769:
			begin
				a25[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			770:
			begin
				a25[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			771:
			begin
				a25[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			772:
			begin
				a25[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			773:
			begin
				a25[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			774:
			begin
				a25[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			775:
			begin
				a25[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			776:
			begin
				a25[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			777:
			begin
				a25[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			778:
			begin
				a25[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			779:
			begin
				a25[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			780:
			begin
				a26[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			781:
			begin
				a26[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			782:
			begin
				a26[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			783:
			begin
				a26[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			784:
			begin
				a26[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			785:
			begin
				a26[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			786:
			begin
				a26[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			787:
			begin
				a26[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			788:
			begin
				a26[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			789:
			begin
				a26[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			790:
			begin
				a26[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			791:
			begin
				a26[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			792:
			begin
				a26[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			793:
			begin
				a26[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			794:
			begin
				a26[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			795:
			begin
				a26[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			796:
			begin
				a26[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			797:
			begin
				a26[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			798:
			begin
				a26[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			799:
			begin
				a26[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			800:
			begin
				a26[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			801:
			begin
				a26[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			802:
			begin
				a26[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			803:
			begin
				a26[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			804:
			begin
				a26[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			805:
			begin
				a26[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			806:
			begin
				a26[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			807:
			begin
				a26[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			808:
			begin
				a26[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			809:
			begin
				a26[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			810:
			begin
				a27[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			811:
			begin
				a27[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			812:
			begin
				a27[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			813:
			begin
				a27[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			814:
			begin
				a27[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			815:
			begin
				a27[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			816:
			begin
				a27[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			817:
			begin
				a27[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			818:
			begin
				a27[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			819:
			begin
				a27[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			820:
			begin
				a27[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			821:
			begin
				a27[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			822:
			begin
				a27[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			823:
			begin
				a27[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			824:
			begin
				a27[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			825:
			begin
				a27[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			826:
			begin
				a27[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			827:
			begin
				a27[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			828:
			begin
				a27[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			829:
			begin
				a27[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			830:
			begin
				a27[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			831:
			begin
				a27[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			832:
			begin
				a27[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			833:
			begin
				a27[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			834:
			begin
				a27[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			835:
			begin
				a27[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			836:
			begin
				a27[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			837:
			begin
				a27[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			838:
			begin
				a27[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			839:
			begin
				a27[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			840:
			begin
				a28[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			841:
			begin
				a28[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			842:
			begin
				a28[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			843:
			begin
				a28[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			844:
			begin
				a28[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			845:
			begin
				a28[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			846:
			begin
				a28[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			847:
			begin
				a28[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			848:
			begin
				a28[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			849:
			begin
				a28[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			850:
			begin
				a28[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			851:
			begin
				a28[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			852:
			begin
				a28[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			853:
			begin
				a28[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			854:
			begin
				a28[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			855:
			begin
				a28[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			856:
			begin
				a28[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			857:
			begin
				a28[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			858:
			begin
				a28[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			859:
			begin
				a28[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			860:
			begin
				a28[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			861:
			begin
				a28[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			862:
			begin
				a28[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			863:
			begin
				a28[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			864:
			begin
				a28[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			865:
			begin
				a28[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			866:
			begin
				a28[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			867:
			begin
				a28[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			868:
			begin
				a28[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			869:
			begin
				a28[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			870:
			begin
				a29[0] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			871:
			begin
				a29[1] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			872:
			begin
				a29[2] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			873:
			begin
				a29[3] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			874:
			begin
				a29[4] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			875:
			begin
				a29[5] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			876:
			begin
				a29[6] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			877:
			begin
				a29[7] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			878:
			begin
				a29[8] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			879:
			begin
				a29[9] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			880:
			begin
				a29[10] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			881:
			begin
				a29[11] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			882:
			begin
				a29[12] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			883:
			begin
				a29[13] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			884:
			begin
				a29[14] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			885:
			begin
				a29[15] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			886:
			begin
				a29[16] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			887:
			begin
				a29[17] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			888:
			begin
				a29[18] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			889:
			begin
				a29[19] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			890:
			begin
				a29[20] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			891:
			begin
				a29[21] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			892:
			begin
				a29[22] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			893:
			begin
				a29[23] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			894:
			begin
				a29[24] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			895:
			begin
				a29[25] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			896:
			begin
				a29[26] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			897:
			begin
				a29[27] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			898:
			begin
				a29[28] <= data_in;
				clk_counter <= clk_counter + 1;
			end
			899:
			begin
				a29[29] <= data_in;
				clk_counter <= clk_counter + 1;
			end
            default: 
        endcase
    end
end

endmodule