`timescale 1ns / 1ps
// memory size 30*30

module mem30x30#(parameter WIDTH = 9)
(
    input clk,
    input rst_n,

    input rd_en,            // read enable
    input wr_en,            // write enable

    input [9:0] rdaddr,     // read address: [9:5] target memline + [4:0] mem address
    input [9:0] wraddr,     // write address: [9:5] target memline + [4:0] mem address

    input [WIDTH-1:0] data_in,

    output [WIDTH-1:0] out
);

// memory
reg [WIDTH-1:0] mem00 [29:0];
reg [WIDTH-1:0] mem01 [29:0];
reg [WIDTH-1:0] mem02 [29:0];
reg [WIDTH-1:0] mem03 [29:0];
reg [WIDTH-1:0] mem04 [29:0];
reg [WIDTH-1:0] mem05 [29:0];
reg [WIDTH-1:0] mem06 [29:0];
reg [WIDTH-1:0] mem07 [29:0];
reg [WIDTH-1:0] mem08 [29:0];
reg [WIDTH-1:0] mem09 [29:0];
reg [WIDTH-1:0] mem10 [29:0];
reg [WIDTH-1:0] mem11 [29:0];
reg [WIDTH-1:0] mem12 [29:0];
reg [WIDTH-1:0] mem13 [29:0];
reg [WIDTH-1:0] mem14 [29:0];
reg [WIDTH-1:0] mem15 [29:0];
reg [WIDTH-1:0] mem16 [29:0];
reg [WIDTH-1:0] mem17 [29:0];
reg [WIDTH-1:0] mem18 [29:0];
reg [WIDTH-1:0] mem19 [29:0];
reg [WIDTH-1:0] mem20 [29:0];
reg [WIDTH-1:0] mem21 [29:0];
reg [WIDTH-1:0] mem22 [29:0];
reg [WIDTH-1:0] mem23 [29:0];
reg [WIDTH-1:0] mem24 [29:0];
reg [WIDTH-1:0] mem25 [29:0];
reg [WIDTH-1:0] mem26 [29:0];
reg [WIDTH-1:0] mem27 [29:0];
reg [WIDTH-1:0] mem28 [29:0];
reg [WIDTH-1:0] mem29 [29:0];

// mem address line
wire [30*WIDTH-1:0] memline00;
wire [30*WIDTH-1:0] memline01;
wire [30*WIDTH-1:0] memline02;
wire [30*WIDTH-1:0] memline03;
wire [30*WIDTH-1:0] memline04;
wire [30*WIDTH-1:0] memline05;
wire [30*WIDTH-1:0] memline06;
wire [30*WIDTH-1:0] memline07;
wire [30*WIDTH-1:0] memline08;
wire [30*WIDTH-1:0] memline09;
wire [30*WIDTH-1:0] memline10;
wire [30*WIDTH-1:0] memline11;
wire [30*WIDTH-1:0] memline12;
wire [30*WIDTH-1:0] memline13;
wire [30*WIDTH-1:0] memline14;
wire [30*WIDTH-1:0] memline15;
wire [30*WIDTH-1:0] memline16;
wire [30*WIDTH-1:0] memline17;
wire [30*WIDTH-1:0] memline18;
wire [30*WIDTH-1:0] memline19;
wire [30*WIDTH-1:0] memline20;
wire [30*WIDTH-1:0] memline21;
wire [30*WIDTH-1:0] memline22;
wire [30*WIDTH-1:0] memline23;
wire [30*WIDTH-1:0] memline24;
wire [30*WIDTH-1:0] memline25;
wire [30*WIDTH-1:0] memline26;
wire [30*WIDTH-1:0] memline27;
wire [30*WIDTH-1:0] memline28;
wire [30*WIDTH-1:0] memline29;

assign memline00 = {mem00[0],mem00[1],mem00[2],mem00[3],mem00[4],mem00[5],mem00[6],mem00[7],mem00[8],mem00[9],mem00[10],mem00[11],mem00[12],mem00[13],mem00[14],mem00[15],mem00[16],mem00[17],mem00[18],mem00[19],mem00[20],mem00[21],mem00[22],mem00[23],mem00[24],mem00[25],mem00[26],mem00[27],mem00[28],mem00[29]};
assign memline01 = {mem01[0],mem01[1],mem01[2],mem01[3],mem01[4],mem01[5],mem01[6],mem01[7],mem01[8],mem01[9],mem01[10],mem01[11],mem01[12],mem01[13],mem01[14],mem01[15],mem01[16],mem01[17],mem01[18],mem01[19],mem01[20],mem01[21],mem01[22],mem01[23],mem01[24],mem01[25],mem01[26],mem01[27],mem01[28],mem01[29]};
assign memline02 = {mem02[0],mem02[1],mem02[2],mem02[3],mem02[4],mem02[5],mem02[6],mem02[7],mem02[8],mem02[9],mem02[10],mem02[11],mem02[12],mem02[13],mem02[14],mem02[15],mem02[16],mem02[17],mem02[18],mem02[19],mem02[20],mem02[21],mem02[22],mem02[23],mem02[24],mem02[25],mem02[26],mem02[27],mem02[28],mem02[29]};
assign memline03 = {mem03[0],mem03[1],mem03[2],mem03[3],mem03[4],mem03[5],mem03[6],mem03[7],mem03[8],mem03[9],mem03[10],mem03[11],mem03[12],mem03[13],mem03[14],mem03[15],mem03[16],mem03[17],mem03[18],mem03[19],mem03[20],mem03[21],mem03[22],mem03[23],mem03[24],mem03[25],mem03[26],mem03[27],mem03[28],mem03[29]};
assign memline04 = {mem04[0],mem04[1],mem04[2],mem04[3],mem04[4],mem04[5],mem04[6],mem04[7],mem04[8],mem04[9],mem04[10],mem04[11],mem04[12],mem04[13],mem04[14],mem04[15],mem04[16],mem04[17],mem04[18],mem04[19],mem04[20],mem04[21],mem04[22],mem04[23],mem04[24],mem04[25],mem04[26],mem04[27],mem04[28],mem04[29]};
assign memline05 = {mem05[0],mem05[1],mem05[2],mem05[3],mem05[4],mem05[5],mem05[6],mem05[7],mem05[8],mem05[9],mem05[10],mem05[11],mem05[12],mem05[13],mem05[14],mem05[15],mem05[16],mem05[17],mem05[18],mem05[19],mem05[20],mem05[21],mem05[22],mem05[23],mem05[24],mem05[25],mem05[26],mem05[27],mem05[28],mem05[29]};
assign memline06 = {mem06[0],mem06[1],mem06[2],mem06[3],mem06[4],mem06[5],mem06[6],mem06[7],mem06[8],mem06[9],mem06[10],mem06[11],mem06[12],mem06[13],mem06[14],mem06[15],mem06[16],mem06[17],mem06[18],mem06[19],mem06[20],mem06[21],mem06[22],mem06[23],mem06[24],mem06[25],mem06[26],mem06[27],mem06[28],mem06[29]};
assign memline07 = {mem07[0],mem07[1],mem07[2],mem07[3],mem07[4],mem07[5],mem07[6],mem07[7],mem07[8],mem07[9],mem07[10],mem07[11],mem07[12],mem07[13],mem07[14],mem07[15],mem07[16],mem07[17],mem07[18],mem07[19],mem07[20],mem07[21],mem07[22],mem07[23],mem07[24],mem07[25],mem07[26],mem07[27],mem07[28],mem07[29]};
assign memline08 = {mem08[0],mem08[1],mem08[2],mem08[3],mem08[4],mem08[5],mem08[6],mem08[7],mem08[8],mem08[9],mem08[10],mem08[11],mem08[12],mem08[13],mem08[14],mem08[15],mem08[16],mem08[17],mem08[18],mem08[19],mem08[20],mem08[21],mem08[22],mem08[23],mem08[24],mem08[25],mem08[26],mem08[27],mem08[28],mem08[29]};
assign memline09 = {mem09[0],mem09[1],mem09[2],mem09[3],mem09[4],mem09[5],mem09[6],mem09[7],mem09[8],mem09[9],mem09[10],mem09[11],mem09[12],mem09[13],mem09[14],mem09[15],mem09[16],mem09[17],mem09[18],mem09[19],mem09[20],mem09[21],mem09[22],mem09[23],mem09[24],mem09[25],mem09[26],mem09[27],mem09[28],mem09[29]};
assign memline10 = {mem10[0],mem10[1],mem10[2],mem10[3],mem10[4],mem10[5],mem10[6],mem10[7],mem10[8],mem10[9],mem10[10],mem10[11],mem10[12],mem10[13],mem10[14],mem10[15],mem10[16],mem10[17],mem10[18],mem10[19],mem10[20],mem10[21],mem10[22],mem10[23],mem10[24],mem10[25],mem10[26],mem10[27],mem10[28],mem10[29]};
assign memline11 = {mem11[0],mem11[1],mem11[2],mem11[3],mem11[4],mem11[5],mem11[6],mem11[7],mem11[8],mem11[9],mem11[10],mem11[11],mem11[12],mem11[13],mem11[14],mem11[15],mem11[16],mem11[17],mem11[18],mem11[19],mem11[20],mem11[21],mem11[22],mem11[23],mem11[24],mem11[25],mem11[26],mem11[27],mem11[28],mem11[29]};
assign memline12 = {mem12[0],mem12[1],mem12[2],mem12[3],mem12[4],mem12[5],mem12[6],mem12[7],mem12[8],mem12[9],mem12[10],mem12[11],mem12[12],mem12[13],mem12[14],mem12[15],mem12[16],mem12[17],mem12[18],mem12[19],mem12[20],mem12[21],mem12[22],mem12[23],mem12[24],mem12[25],mem12[26],mem12[27],mem12[28],mem12[29]};
assign memline13 = {mem13[0],mem13[1],mem13[2],mem13[3],mem13[4],mem13[5],mem13[6],mem13[7],mem13[8],mem13[9],mem13[10],mem13[11],mem13[12],mem13[13],mem13[14],mem13[15],mem13[16],mem13[17],mem13[18],mem13[19],mem13[20],mem13[21],mem13[22],mem13[23],mem13[24],mem13[25],mem13[26],mem13[27],mem13[28],mem13[29]};
assign memline14 = {mem14[0],mem14[1],mem14[2],mem14[3],mem14[4],mem14[5],mem14[6],mem14[7],mem14[8],mem14[9],mem14[10],mem14[11],mem14[12],mem14[13],mem14[14],mem14[15],mem14[16],mem14[17],mem14[18],mem14[19],mem14[20],mem14[21],mem14[22],mem14[23],mem14[24],mem14[25],mem14[26],mem14[27],mem14[28],mem14[29]};
assign memline15 = {mem15[0],mem15[1],mem15[2],mem15[3],mem15[4],mem15[5],mem15[6],mem15[7],mem15[8],mem15[9],mem15[10],mem15[11],mem15[12],mem15[13],mem15[14],mem15[15],mem15[16],mem15[17],mem15[18],mem15[19],mem15[20],mem15[21],mem15[22],mem15[23],mem15[24],mem15[25],mem15[26],mem15[27],mem15[28],mem15[29]};
assign memline16 = {mem16[0],mem16[1],mem16[2],mem16[3],mem16[4],mem16[5],mem16[6],mem16[7],mem16[8],mem16[9],mem16[10],mem16[11],mem16[12],mem16[13],mem16[14],mem16[15],mem16[16],mem16[17],mem16[18],mem16[19],mem16[20],mem16[21],mem16[22],mem16[23],mem16[24],mem16[25],mem16[26],mem16[27],mem16[28],mem16[29]};
assign memline17 = {mem17[0],mem17[1],mem17[2],mem17[3],mem17[4],mem17[5],mem17[6],mem17[7],mem17[8],mem17[9],mem17[10],mem17[11],mem17[12],mem17[13],mem17[14],mem17[15],mem17[16],mem17[17],mem17[18],mem17[19],mem17[20],mem17[21],mem17[22],mem17[23],mem17[24],mem17[25],mem17[26],mem17[27],mem17[28],mem17[29]};
assign memline18 = {mem18[0],mem18[1],mem18[2],mem18[3],mem18[4],mem18[5],mem18[6],mem18[7],mem18[8],mem18[9],mem18[10],mem18[11],mem18[12],mem18[13],mem18[14],mem18[15],mem18[16],mem18[17],mem18[18],mem18[19],mem18[20],mem18[21],mem18[22],mem18[23],mem18[24],mem18[25],mem18[26],mem18[27],mem18[28],mem18[29]};
assign memline19 = {mem19[0],mem19[1],mem19[2],mem19[3],mem19[4],mem19[5],mem19[6],mem19[7],mem19[8],mem19[9],mem19[10],mem19[11],mem19[12],mem19[13],mem19[14],mem19[15],mem19[16],mem19[17],mem19[18],mem19[19],mem19[20],mem19[21],mem19[22],mem19[23],mem19[24],mem19[25],mem19[26],mem19[27],mem19[28],mem19[29]};
assign memline20 = {mem20[0],mem20[1],mem20[2],mem20[3],mem20[4],mem20[5],mem20[6],mem20[7],mem20[8],mem20[9],mem20[10],mem20[11],mem20[12],mem20[13],mem20[14],mem20[15],mem20[16],mem20[17],mem20[18],mem20[19],mem20[20],mem20[21],mem20[22],mem20[23],mem20[24],mem20[25],mem20[26],mem20[27],mem20[28],mem20[29]};
assign memline21 = {mem21[0],mem21[1],mem21[2],mem21[3],mem21[4],mem21[5],mem21[6],mem21[7],mem21[8],mem21[9],mem21[10],mem21[11],mem21[12],mem21[13],mem21[14],mem21[15],mem21[16],mem21[17],mem21[18],mem21[19],mem21[20],mem21[21],mem21[22],mem21[23],mem21[24],mem21[25],mem21[26],mem21[27],mem21[28],mem21[29]};
assign memline22 = {mem22[0],mem22[1],mem22[2],mem22[3],mem22[4],mem22[5],mem22[6],mem22[7],mem22[8],mem22[9],mem22[10],mem22[11],mem22[12],mem22[13],mem22[14],mem22[15],mem22[16],mem22[17],mem22[18],mem22[19],mem22[20],mem22[21],mem22[22],mem22[23],mem22[24],mem22[25],mem22[26],mem22[27],mem22[28],mem22[29]};
assign memline23 = {mem23[0],mem23[1],mem23[2],mem23[3],mem23[4],mem23[5],mem23[6],mem23[7],mem23[8],mem23[9],mem23[10],mem23[11],mem23[12],mem23[13],mem23[14],mem23[15],mem23[16],mem23[17],mem23[18],mem23[19],mem23[20],mem23[21],mem23[22],mem23[23],mem23[24],mem23[25],mem23[26],mem23[27],mem23[28],mem23[29]};
assign memline24 = {mem24[0],mem24[1],mem24[2],mem24[3],mem24[4],mem24[5],mem24[6],mem24[7],mem24[8],mem24[9],mem24[10],mem24[11],mem24[12],mem24[13],mem24[14],mem24[15],mem24[16],mem24[17],mem24[18],mem24[19],mem24[20],mem24[21],mem24[22],mem24[23],mem24[24],mem24[25],mem24[26],mem24[27],mem24[28],mem24[29]};
assign memline25 = {mem25[0],mem25[1],mem25[2],mem25[3],mem25[4],mem25[5],mem25[6],mem25[7],mem25[8],mem25[9],mem25[10],mem25[11],mem25[12],mem25[13],mem25[14],mem25[15],mem25[16],mem25[17],mem25[18],mem25[19],mem25[20],mem25[21],mem25[22],mem25[23],mem25[24],mem25[25],mem25[26],mem25[27],mem25[28],mem25[29]};
assign memline26 = {mem26[0],mem26[1],mem26[2],mem26[3],mem26[4],mem26[5],mem26[6],mem26[7],mem26[8],mem26[9],mem26[10],mem26[11],mem26[12],mem26[13],mem26[14],mem26[15],mem26[16],mem26[17],mem26[18],mem26[19],mem26[20],mem26[21],mem26[22],mem26[23],mem26[24],mem26[25],mem26[26],mem26[27],mem26[28],mem26[29]};
assign memline27 = {mem27[0],mem27[1],mem27[2],mem27[3],mem27[4],mem27[5],mem27[6],mem27[7],mem27[8],mem27[9],mem27[10],mem27[11],mem27[12],mem27[13],mem27[14],mem27[15],mem27[16],mem27[17],mem27[18],mem27[19],mem27[20],mem27[21],mem27[22],mem27[23],mem27[24],mem27[25],mem27[26],mem27[27],mem27[28],mem27[29]};
assign memline28 = {mem28[0],mem28[1],mem28[2],mem28[3],mem28[4],mem28[5],mem28[6],mem28[7],mem28[8],mem28[9],mem28[10],mem28[11],mem28[12],mem28[13],mem28[14],mem28[15],mem28[16],mem28[17],mem28[18],mem28[19],mem28[20],mem28[21],mem28[22],mem28[23],mem28[24],mem28[25],mem28[26],mem28[27],mem28[28],mem28[29]};
assign memline29 = {mem29[0],mem29[1],mem29[2],mem29[3],mem29[4],mem29[5],mem29[6],mem29[7],mem29[8],mem29[9],mem29[10],mem29[11],mem29[12],mem29[13],mem29[14],mem29[15],mem29[16],mem29[17],mem29[18],mem29[19],mem29[20],mem29[21],mem29[22],mem29[23],mem29[24],mem29[25],mem29[26],mem29[27],mem29[28],mem29[29]};



/**********************************************************************************************************************/
/************************************************ READ & WRITE Logic **************************************************/
/**********************************************************************************************************************/
reg [4:0] target_line;
reg [4:0] addr;
reg [WIDTH-1:0] out_buffer;

initial
begin
    target_line = 5'b00000;
    addr = 5'b00000;
end

// resolve target line
always@(posedge clk)
begin
    if(rd_en) begin
        target_line <= rdaddr[9:5];
        addr <= rdaddr[4:0];
    end
    else if(wr_en) begin
        target_line <= wraddr[9:5];
        addr <= wraddr[4:0];
    end
    else begin
        target_line <= 5'b00000;
        addr <= 5'b00000;
    end
end

always@(posedge clk or negedge rst_n)
begin
    if(rst_n)
        out_buffer <= 0;
    else if(rd_en)
        case (target_line)
			0:
			case(addr)
				0:out_buffer <= mem00[0];
				1:out_buffer <= mem00[1];
				2:out_buffer <= mem00[2];
				3:out_buffer <= mem00[3];
				4:out_buffer <= mem00[4];
				5:out_buffer <= mem00[5];
				6:out_buffer <= mem00[6];
				7:out_buffer <= mem00[7];
				8:out_buffer <= mem00[8];
				9:out_buffer <= mem00[9];
				10:out_buffer <= mem00[10];
				11:out_buffer <= mem00[11];
				12:out_buffer <= mem00[12];
				13:out_buffer <= mem00[13];
				14:out_buffer <= mem00[14];
				15:out_buffer <= mem00[15];
				16:out_buffer <= mem00[16];
				17:out_buffer <= mem00[17];
				18:out_buffer <= mem00[18];
				19:out_buffer <= mem00[19];
				20:out_buffer <= mem00[20];
				21:out_buffer <= mem00[21];
				22:out_buffer <= mem00[22];
				23:out_buffer <= mem00[23];
				24:out_buffer <= mem00[24];
				25:out_buffer <= mem00[25];
				26:out_buffer <= mem00[26];
				27:out_buffer <= mem00[27];
				28:out_buffer <= mem00[28];
				29:out_buffer <= mem00[29];
			endcase
		
			1:
			case(addr)
				0:out_buffer <= mem01[0];
				1:out_buffer <= mem01[1];
				2:out_buffer <= mem01[2];
				3:out_buffer <= mem01[3];
				4:out_buffer <= mem01[4];
				5:out_buffer <= mem01[5];
				6:out_buffer <= mem01[6];
				7:out_buffer <= mem01[7];
				8:out_buffer <= mem01[8];
				9:out_buffer <= mem01[9];
				10:out_buffer <= mem01[10];
				11:out_buffer <= mem01[11];
				12:out_buffer <= mem01[12];
				13:out_buffer <= mem01[13];
				14:out_buffer <= mem01[14];
				15:out_buffer <= mem01[15];
				16:out_buffer <= mem01[16];
				17:out_buffer <= mem01[17];
				18:out_buffer <= mem01[18];
				19:out_buffer <= mem01[19];
				20:out_buffer <= mem01[20];
				21:out_buffer <= mem01[21];
				22:out_buffer <= mem01[22];
				23:out_buffer <= mem01[23];
				24:out_buffer <= mem01[24];
				25:out_buffer <= mem01[25];
				26:out_buffer <= mem01[26];
				27:out_buffer <= mem01[27];
				28:out_buffer <= mem01[28];
				29:out_buffer <= mem01[29];
			endcase
		
			2:
			case(addr)
				0:out_buffer <= mem02[0];
				1:out_buffer <= mem02[1];
				2:out_buffer <= mem02[2];
				3:out_buffer <= mem02[3];
				4:out_buffer <= mem02[4];
				5:out_buffer <= mem02[5];
				6:out_buffer <= mem02[6];
				7:out_buffer <= mem02[7];
				8:out_buffer <= mem02[8];
				9:out_buffer <= mem02[9];
				10:out_buffer <= mem02[10];
				11:out_buffer <= mem02[11];
				12:out_buffer <= mem02[12];
				13:out_buffer <= mem02[13];
				14:out_buffer <= mem02[14];
				15:out_buffer <= mem02[15];
				16:out_buffer <= mem02[16];
				17:out_buffer <= mem02[17];
				18:out_buffer <= mem02[18];
				19:out_buffer <= mem02[19];
				20:out_buffer <= mem02[20];
				21:out_buffer <= mem02[21];
				22:out_buffer <= mem02[22];
				23:out_buffer <= mem02[23];
				24:out_buffer <= mem02[24];
				25:out_buffer <= mem02[25];
				26:out_buffer <= mem02[26];
				27:out_buffer <= mem02[27];
				28:out_buffer <= mem02[28];
				29:out_buffer <= mem02[29];
			endcase
			
			3:
			case(addr)
				0:out_buffer <= mem03[0];
				1:out_buffer <= mem03[1];
				2:out_buffer <= mem03[2];
				3:out_buffer <= mem03[3];
				4:out_buffer <= mem03[4];
				5:out_buffer <= mem03[5];
				6:out_buffer <= mem03[6];
				7:out_buffer <= mem03[7];
				8:out_buffer <= mem03[8];
				9:out_buffer <= mem03[9];
				10:out_buffer <= mem03[10];
				11:out_buffer <= mem03[11];
				12:out_buffer <= mem03[12];
				13:out_buffer <= mem03[13];
				14:out_buffer <= mem03[14];
				15:out_buffer <= mem03[15];
				16:out_buffer <= mem03[16];
				17:out_buffer <= mem03[17];
				18:out_buffer <= mem03[18];
				19:out_buffer <= mem03[19];
				20:out_buffer <= mem03[20];
				21:out_buffer <= mem03[21];
				22:out_buffer <= mem03[22];
				23:out_buffer <= mem03[23];
				24:out_buffer <= mem03[24];
				25:out_buffer <= mem03[25];
				26:out_buffer <= mem03[26];
				27:out_buffer <= mem03[27];
				28:out_buffer <= mem03[28];
				29:out_buffer <= mem03[29];
			endcase
			
			4:
			case(addr)
				0:out_buffer <= mem04[0];
				1:out_buffer <= mem04[1];
				2:out_buffer <= mem04[2];
				3:out_buffer <= mem04[3];
				4:out_buffer <= mem04[4];
				5:out_buffer <= mem04[5];
				6:out_buffer <= mem04[6];
				7:out_buffer <= mem04[7];
				8:out_buffer <= mem04[8];
				9:out_buffer <= mem04[9];
				10:out_buffer <= mem04[10];
				11:out_buffer <= mem04[11];
				12:out_buffer <= mem04[12];
				13:out_buffer <= mem04[13];
				14:out_buffer <= mem04[14];
				15:out_buffer <= mem04[15];
				16:out_buffer <= mem04[16];
				17:out_buffer <= mem04[17];
				18:out_buffer <= mem04[18];
				19:out_buffer <= mem04[19];
				20:out_buffer <= mem04[20];
				21:out_buffer <= mem04[21];
				22:out_buffer <= mem04[22];
				23:out_buffer <= mem04[23];
				24:out_buffer <= mem04[24];
				25:out_buffer <= mem04[25];
				26:out_buffer <= mem04[26];
				27:out_buffer <= mem04[27];
				28:out_buffer <= mem04[28];
				29:out_buffer <= mem04[29];
			endcase
			
			5:
			case(addr)
				0:out_buffer <= mem05[0];
				1:out_buffer <= mem05[1];
				2:out_buffer <= mem05[2];
				3:out_buffer <= mem05[3];
				4:out_buffer <= mem05[4];
				5:out_buffer <= mem05[5];
				6:out_buffer <= mem05[6];
				7:out_buffer <= mem05[7];
				8:out_buffer <= mem05[8];
				9:out_buffer <= mem05[9];
				10:out_buffer <= mem05[10];
				11:out_buffer <= mem05[11];
				12:out_buffer <= mem05[12];
				13:out_buffer <= mem05[13];
				14:out_buffer <= mem05[14];
				15:out_buffer <= mem05[15];
				16:out_buffer <= mem05[16];
				17:out_buffer <= mem05[17];
				18:out_buffer <= mem05[18];
				19:out_buffer <= mem05[19];
				20:out_buffer <= mem05[20];
				21:out_buffer <= mem05[21];
				22:out_buffer <= mem05[22];
				23:out_buffer <= mem05[23];
				24:out_buffer <= mem05[24];
				25:out_buffer <= mem05[25];
				26:out_buffer <= mem05[26];
				27:out_buffer <= mem05[27];
				28:out_buffer <= mem05[28];
				29:out_buffer <= mem05[29];
			endcase
			
			6:
			case(addr)
				0:out_buffer <= mem06[0];
				1:out_buffer <= mem06[1];
				2:out_buffer <= mem06[2];
				3:out_buffer <= mem06[3];
				4:out_buffer <= mem06[4];
				5:out_buffer <= mem06[5];
				6:out_buffer <= mem06[6];
				7:out_buffer <= mem06[7];
				8:out_buffer <= mem06[8];
				9:out_buffer <= mem06[9];
				10:out_buffer <= mem06[10];
				11:out_buffer <= mem06[11];
				12:out_buffer <= mem06[12];
				13:out_buffer <= mem06[13];
				14:out_buffer <= mem06[14];
				15:out_buffer <= mem06[15];
				16:out_buffer <= mem06[16];
				17:out_buffer <= mem06[17];
				18:out_buffer <= mem06[18];
				19:out_buffer <= mem06[19];
				20:out_buffer <= mem06[20];
				21:out_buffer <= mem06[21];
				22:out_buffer <= mem06[22];
				23:out_buffer <= mem06[23];
				24:out_buffer <= mem06[24];
				25:out_buffer <= mem06[25];
				26:out_buffer <= mem06[26];
				27:out_buffer <= mem06[27];
				28:out_buffer <= mem06[28];
				29:out_buffer <= mem06[29];
			endcase
			
			7:
			case(addr)
				0:out_buffer <= mem07[0];
				1:out_buffer <= mem07[1];
				2:out_buffer <= mem07[2];
				3:out_buffer <= mem07[3];
				4:out_buffer <= mem07[4];
				5:out_buffer <= mem07[5];
				6:out_buffer <= mem07[6];
				7:out_buffer <= mem07[7];
				8:out_buffer <= mem07[8];
				9:out_buffer <= mem07[9];
				10:out_buffer <= mem07[10];
				11:out_buffer <= mem07[11];
				12:out_buffer <= mem07[12];
				13:out_buffer <= mem07[13];
				14:out_buffer <= mem07[14];
				15:out_buffer <= mem07[15];
				16:out_buffer <= mem07[16];
				17:out_buffer <= mem07[17];
				18:out_buffer <= mem07[18];
				19:out_buffer <= mem07[19];
				20:out_buffer <= mem07[20];
				21:out_buffer <= mem07[21];
				22:out_buffer <= mem07[22];
				23:out_buffer <= mem07[23];
				24:out_buffer <= mem07[24];
				25:out_buffer <= mem07[25];
				26:out_buffer <= mem07[26];
				27:out_buffer <= mem07[27];
				28:out_buffer <= mem07[28];
				29:out_buffer <= mem07[29];
			endcase
			
			8:
			case(addr)
				0:out_buffer <= mem08[0];
				1:out_buffer <= mem08[1];
				2:out_buffer <= mem08[2];
				3:out_buffer <= mem08[3];
				4:out_buffer <= mem08[4];
				5:out_buffer <= mem08[5];
				6:out_buffer <= mem08[6];
				7:out_buffer <= mem08[7];
				8:out_buffer <= mem08[8];
				9:out_buffer <= mem08[9];
				10:out_buffer <= mem08[10];
				11:out_buffer <= mem08[11];
				12:out_buffer <= mem08[12];
				13:out_buffer <= mem08[13];
				14:out_buffer <= mem08[14];
				15:out_buffer <= mem08[15];
				16:out_buffer <= mem08[16];
				17:out_buffer <= mem08[17];
				18:out_buffer <= mem08[18];
				19:out_buffer <= mem08[19];
				20:out_buffer <= mem08[20];
				21:out_buffer <= mem08[21];
				22:out_buffer <= mem08[22];
				23:out_buffer <= mem08[23];
				24:out_buffer <= mem08[24];
				25:out_buffer <= mem08[25];
				26:out_buffer <= mem08[26];
				27:out_buffer <= mem08[27];
				28:out_buffer <= mem08[28];
				29:out_buffer <= mem08[29];
			endcase
			
			9:
			case(addr)
				0:out_buffer <= mem09[0];
				1:out_buffer <= mem09[1];
				2:out_buffer <= mem09[2];
				3:out_buffer <= mem09[3];
				4:out_buffer <= mem09[4];
				5:out_buffer <= mem09[5];
				6:out_buffer <= mem09[6];
				7:out_buffer <= mem09[7];
				8:out_buffer <= mem09[8];
				9:out_buffer <= mem09[9];
				10:out_buffer <= mem09[10];
				11:out_buffer <= mem09[11];
				12:out_buffer <= mem09[12];
				13:out_buffer <= mem09[13];
				14:out_buffer <= mem09[14];
				15:out_buffer <= mem09[15];
				16:out_buffer <= mem09[16];
				17:out_buffer <= mem09[17];
				18:out_buffer <= mem09[18];
				19:out_buffer <= mem09[19];
				20:out_buffer <= mem09[20];
				21:out_buffer <= mem09[21];
				22:out_buffer <= mem09[22];
				23:out_buffer <= mem09[23];
				24:out_buffer <= mem09[24];
				25:out_buffer <= mem09[25];
				26:out_buffer <= mem09[26];
				27:out_buffer <= mem09[27];
				28:out_buffer <= mem09[28];
				29:out_buffer <= mem09[29];
			endcase
			
			10:
			case(addr)
				0:out_buffer <= mem10[0];
				1:out_buffer <= mem10[1];
				2:out_buffer <= mem10[2];
				3:out_buffer <= mem10[3];
				4:out_buffer <= mem10[4];
				5:out_buffer <= mem10[5];
				6:out_buffer <= mem10[6];
				7:out_buffer <= mem10[7];
				8:out_buffer <= mem10[8];
				9:out_buffer <= mem10[9];
				10:out_buffer <= mem10[10];
				11:out_buffer <= mem10[11];
				12:out_buffer <= mem10[12];
				13:out_buffer <= mem10[13];
				14:out_buffer <= mem10[14];
				15:out_buffer <= mem10[15];
				16:out_buffer <= mem10[16];
				17:out_buffer <= mem10[17];
				18:out_buffer <= mem10[18];
				19:out_buffer <= mem10[19];
				20:out_buffer <= mem10[20];
				21:out_buffer <= mem10[21];
				22:out_buffer <= mem10[22];
				23:out_buffer <= mem10[23];
				24:out_buffer <= mem10[24];
				25:out_buffer <= mem10[25];
				26:out_buffer <= mem10[26];
				27:out_buffer <= mem10[27];
				28:out_buffer <= mem10[28];
				29:out_buffer <= mem10[29];
			endcase
			
			11:
			case(addr)
				0:out_buffer <= mem11[0];
				1:out_buffer <= mem11[1];
				2:out_buffer <= mem11[2];
				3:out_buffer <= mem11[3];
				4:out_buffer <= mem11[4];
				5:out_buffer <= mem11[5];
				6:out_buffer <= mem11[6];
				7:out_buffer <= mem11[7];
				8:out_buffer <= mem11[8];
				9:out_buffer <= mem11[9];
				10:out_buffer <= mem11[10];
				11:out_buffer <= mem11[11];
				12:out_buffer <= mem11[12];
				13:out_buffer <= mem11[13];
				14:out_buffer <= mem11[14];
				15:out_buffer <= mem11[15];
				16:out_buffer <= mem11[16];
				17:out_buffer <= mem11[17];
				18:out_buffer <= mem11[18];
				19:out_buffer <= mem11[19];
				20:out_buffer <= mem11[20];
				21:out_buffer <= mem11[21];
				22:out_buffer <= mem11[22];
				23:out_buffer <= mem11[23];
				24:out_buffer <= mem11[24];
				25:out_buffer <= mem11[25];
				26:out_buffer <= mem11[26];
				27:out_buffer <= mem11[27];
				28:out_buffer <= mem11[28];
				29:out_buffer <= mem11[29];
			endcase

			12:
			case(addr)
				0:out_buffer <= mem12[0];
				1:out_buffer <= mem12[1];
				2:out_buffer <= mem12[2];
				3:out_buffer <= mem12[3];
				4:out_buffer <= mem12[4];
				5:out_buffer <= mem12[5];
				6:out_buffer <= mem12[6];
				7:out_buffer <= mem12[7];
				8:out_buffer <= mem12[8];
				9:out_buffer <= mem12[9];
				10:out_buffer <= mem12[10];
				11:out_buffer <= mem12[11];
				12:out_buffer <= mem12[12];
				13:out_buffer <= mem12[13];
				14:out_buffer <= mem12[14];
				15:out_buffer <= mem12[15];
				16:out_buffer <= mem12[16];
				17:out_buffer <= mem12[17];
				18:out_buffer <= mem12[18];
				19:out_buffer <= mem12[19];
				20:out_buffer <= mem12[20];
				21:out_buffer <= mem12[21];
				22:out_buffer <= mem12[22];
				23:out_buffer <= mem12[23];
				24:out_buffer <= mem12[24];
				25:out_buffer <= mem12[25];
				26:out_buffer <= mem12[26];
				27:out_buffer <= mem12[27];
				28:out_buffer <= mem12[28];
				29:out_buffer <= mem12[29];
			endcase

			13:
			case(addr)
				0:out_buffer <= mem13[0];
				1:out_buffer <= mem13[1];
				2:out_buffer <= mem13[2];
				3:out_buffer <= mem13[3];
				4:out_buffer <= mem13[4];
				5:out_buffer <= mem13[5];
				6:out_buffer <= mem13[6];
				7:out_buffer <= mem13[7];
				8:out_buffer <= mem13[8];
				9:out_buffer <= mem13[9];
				10:out_buffer <= mem13[10];
				11:out_buffer <= mem13[11];
				12:out_buffer <= mem13[12];
				13:out_buffer <= mem13[13];
				14:out_buffer <= mem13[14];
				15:out_buffer <= mem13[15];
				16:out_buffer <= mem13[16];
				17:out_buffer <= mem13[17];
				18:out_buffer <= mem13[18];
				19:out_buffer <= mem13[19];
				20:out_buffer <= mem13[20];
				21:out_buffer <= mem13[21];
				22:out_buffer <= mem13[22];
				23:out_buffer <= mem13[23];
				24:out_buffer <= mem13[24];
				25:out_buffer <= mem13[25];
				26:out_buffer <= mem13[26];
				27:out_buffer <= mem13[27];
				28:out_buffer <= mem13[28];
				29:out_buffer <= mem13[29];
			endcase
			
			14:
			case(addr)
				0:out_buffer <= mem14[0];
				1:out_buffer <= mem14[1];
				2:out_buffer <= mem14[2];
				3:out_buffer <= mem14[3];
				4:out_buffer <= mem14[4];
				5:out_buffer <= mem14[5];
				6:out_buffer <= mem14[6];
				7:out_buffer <= mem14[7];
				8:out_buffer <= mem14[8];
				9:out_buffer <= mem14[9];
				10:out_buffer <= mem14[10];
				11:out_buffer <= mem14[11];
				12:out_buffer <= mem14[12];
				13:out_buffer <= mem14[13];
				14:out_buffer <= mem14[14];
				15:out_buffer <= mem14[15];
				16:out_buffer <= mem14[16];
				17:out_buffer <= mem14[17];
				18:out_buffer <= mem14[18];
				19:out_buffer <= mem14[19];
				20:out_buffer <= mem14[20];
				21:out_buffer <= mem14[21];
				22:out_buffer <= mem14[22];
				23:out_buffer <= mem14[23];
				24:out_buffer <= mem14[24];
				25:out_buffer <= mem14[25];
				26:out_buffer <= mem14[26];
				27:out_buffer <= mem14[27];
				28:out_buffer <= mem14[28];
				29:out_buffer <= mem14[29];
			endcase
			
			15:
			case(addr)
				0:out_buffer <= mem15[0];
				1:out_buffer <= mem15[1];
				2:out_buffer <= mem15[2];
				3:out_buffer <= mem15[3];
				4:out_buffer <= mem15[4];
				5:out_buffer <= mem15[5];
				6:out_buffer <= mem15[6];
				7:out_buffer <= mem15[7];
				8:out_buffer <= mem15[8];
				9:out_buffer <= mem15[9];
				10:out_buffer <= mem15[10];
				11:out_buffer <= mem15[11];
				12:out_buffer <= mem15[12];
				13:out_buffer <= mem15[13];
				14:out_buffer <= mem15[14];
				15:out_buffer <= mem15[15];
				16:out_buffer <= mem15[16];
				17:out_buffer <= mem15[17];
				18:out_buffer <= mem15[18];
				19:out_buffer <= mem15[19];
				20:out_buffer <= mem15[20];
				21:out_buffer <= mem15[21];
				22:out_buffer <= mem15[22];
				23:out_buffer <= mem15[23];
				24:out_buffer <= mem15[24];
				25:out_buffer <= mem15[25];
				26:out_buffer <= mem15[26];
				27:out_buffer <= mem15[27];
				28:out_buffer <= mem15[28];
				29:out_buffer <= mem15[29];
			endcase
			
			16:
			case(addr)
				0:out_buffer <= mem16[0];
				1:out_buffer <= mem16[1];
				2:out_buffer <= mem16[2];
				3:out_buffer <= mem16[3];
				4:out_buffer <= mem16[4];
				5:out_buffer <= mem16[5];
				6:out_buffer <= mem16[6];
				7:out_buffer <= mem16[7];
				8:out_buffer <= mem16[8];
				9:out_buffer <= mem16[9];
				10:out_buffer <= mem16[10];
				11:out_buffer <= mem16[11];
				12:out_buffer <= mem16[12];
				13:out_buffer <= mem16[13];
				14:out_buffer <= mem16[14];
				15:out_buffer <= mem16[15];
				16:out_buffer <= mem16[16];
				17:out_buffer <= mem16[17];
				18:out_buffer <= mem16[18];
				19:out_buffer <= mem16[19];
				20:out_buffer <= mem16[20];
				21:out_buffer <= mem16[21];
				22:out_buffer <= mem16[22];
				23:out_buffer <= mem16[23];
				24:out_buffer <= mem16[24];
				25:out_buffer <= mem16[25];
				26:out_buffer <= mem16[26];
				27:out_buffer <= mem16[27];
				28:out_buffer <= mem16[28];
				29:out_buffer <= mem16[29];
			endcase
		
			17:
			case(addr)
				0:out_buffer <= mem17[0];
				1:out_buffer <= mem17[1];
				2:out_buffer <= mem17[2];
				3:out_buffer <= mem17[3];
				4:out_buffer <= mem17[4];
				5:out_buffer <= mem17[5];
				6:out_buffer <= mem17[6];
				7:out_buffer <= mem17[7];
				8:out_buffer <= mem17[8];
				9:out_buffer <= mem17[9];
				10:out_buffer <= mem17[10];
				11:out_buffer <= mem17[11];
				12:out_buffer <= mem17[12];
				13:out_buffer <= mem17[13];
				14:out_buffer <= mem17[14];
				15:out_buffer <= mem17[15];
				16:out_buffer <= mem17[16];
				17:out_buffer <= mem17[17];
				18:out_buffer <= mem17[18];
				19:out_buffer <= mem17[19];
				20:out_buffer <= mem17[20];
				21:out_buffer <= mem17[21];
				22:out_buffer <= mem17[22];
				23:out_buffer <= mem17[23];
				24:out_buffer <= mem17[24];
				25:out_buffer <= mem17[25];
				26:out_buffer <= mem17[26];
				27:out_buffer <= mem17[27];
				28:out_buffer <= mem17[28];
				29:out_buffer <= mem17[29];
			endcase
		
			18:
			case(addr)
				0:out_buffer <= mem18[0];
				1:out_buffer <= mem18[1];
				2:out_buffer <= mem18[2];
				3:out_buffer <= mem18[3];
				4:out_buffer <= mem18[4];
				5:out_buffer <= mem18[5];
				6:out_buffer <= mem18[6];
				7:out_buffer <= mem18[7];
				8:out_buffer <= mem18[8];
				9:out_buffer <= mem18[9];
				10:out_buffer <= mem18[10];
				11:out_buffer <= mem18[11];
				12:out_buffer <= mem18[12];
				13:out_buffer <= mem18[13];
				14:out_buffer <= mem18[14];
				15:out_buffer <= mem18[15];
				16:out_buffer <= mem18[16];
				17:out_buffer <= mem18[17];
				18:out_buffer <= mem18[18];
				19:out_buffer <= mem18[19];
				20:out_buffer <= mem18[20];
				21:out_buffer <= mem18[21];
				22:out_buffer <= mem18[22];
				23:out_buffer <= mem18[23];
				24:out_buffer <= mem18[24];
				25:out_buffer <= mem18[25];
				26:out_buffer <= mem18[26];
				27:out_buffer <= mem18[27];
				28:out_buffer <= mem18[28];
				29:out_buffer <= mem18[29];
			endcase
		
			19:
			case(addr)
				0:out_buffer <= mem19[0];
				1:out_buffer <= mem19[1];
				2:out_buffer <= mem19[2];
				3:out_buffer <= mem19[3];
				4:out_buffer <= mem19[4];
				5:out_buffer <= mem19[5];
				6:out_buffer <= mem19[6];
				7:out_buffer <= mem19[7];
				8:out_buffer <= mem19[8];
				9:out_buffer <= mem19[9];
				10:out_buffer <= mem19[10];
				11:out_buffer <= mem19[11];
				12:out_buffer <= mem19[12];
				13:out_buffer <= mem19[13];
				14:out_buffer <= mem19[14];
				15:out_buffer <= mem19[15];
				16:out_buffer <= mem19[16];
				17:out_buffer <= mem19[17];
				18:out_buffer <= mem19[18];
				19:out_buffer <= mem19[19];
				20:out_buffer <= mem19[20];
				21:out_buffer <= mem19[21];
				22:out_buffer <= mem19[22];
				23:out_buffer <= mem19[23];
				24:out_buffer <= mem19[24];
				25:out_buffer <= mem19[25];
				26:out_buffer <= mem19[26];
				27:out_buffer <= mem19[27];
				28:out_buffer <= mem19[28];
				29:out_buffer <= mem19[29];
			endcase
			
			20:
			case(addr)
				0:out_buffer <= mem20[0];
				1:out_buffer <= mem20[1];
				2:out_buffer <= mem20[2];
				3:out_buffer <= mem20[3];
				4:out_buffer <= mem20[4];
				5:out_buffer <= mem20[5];
				6:out_buffer <= mem20[6];
				7:out_buffer <= mem20[7];
				8:out_buffer <= mem20[8];
				9:out_buffer <= mem20[9];
				10:out_buffer <= mem20[10];
				11:out_buffer <= mem20[11];
				12:out_buffer <= mem20[12];
				13:out_buffer <= mem20[13];
				14:out_buffer <= mem20[14];
				15:out_buffer <= mem20[15];
				16:out_buffer <= mem20[16];
				17:out_buffer <= mem20[17];
				18:out_buffer <= mem20[18];
				19:out_buffer <= mem20[19];
				20:out_buffer <= mem20[20];
				21:out_buffer <= mem20[21];
				22:out_buffer <= mem20[22];
				23:out_buffer <= mem20[23];
				24:out_buffer <= mem20[24];
				25:out_buffer <= mem20[25];
				26:out_buffer <= mem20[26];
				27:out_buffer <= mem20[27];
				28:out_buffer <= mem20[28];
				29:out_buffer <= mem20[29];
			endcase
		
			21:
			case(addr)
				0:out_buffer <= mem21[0];
				1:out_buffer <= mem21[1];
				2:out_buffer <= mem21[2];
				3:out_buffer <= mem21[3];
				4:out_buffer <= mem21[4];
				5:out_buffer <= mem21[5];
				6:out_buffer <= mem21[6];
				7:out_buffer <= mem21[7];
				8:out_buffer <= mem21[8];
				9:out_buffer <= mem21[9];
				10:out_buffer <= mem21[10];
				11:out_buffer <= mem21[11];
				12:out_buffer <= mem21[12];
				13:out_buffer <= mem21[13];
				14:out_buffer <= mem21[14];
				15:out_buffer <= mem21[15];
				16:out_buffer <= mem21[16];
				17:out_buffer <= mem21[17];
				18:out_buffer <= mem21[18];
				19:out_buffer <= mem21[19];
				20:out_buffer <= mem21[20];
				21:out_buffer <= mem21[21];
				22:out_buffer <= mem21[22];
				23:out_buffer <= mem21[23];
				24:out_buffer <= mem21[24];
				25:out_buffer <= mem21[25];
				26:out_buffer <= mem21[26];
				27:out_buffer <= mem21[27];
				28:out_buffer <= mem21[28];
				29:out_buffer <= mem21[29];
			endcase
		
			22:
			case(addr)
				0:out_buffer <= mem22[0];
				1:out_buffer <= mem22[1];
				2:out_buffer <= mem22[2];
				3:out_buffer <= mem22[3];
				4:out_buffer <= mem22[4];
				5:out_buffer <= mem22[5];
				6:out_buffer <= mem22[6];
				7:out_buffer <= mem22[7];
				8:out_buffer <= mem22[8];
				9:out_buffer <= mem22[9];
				10:out_buffer <= mem22[10];
				11:out_buffer <= mem22[11];
				12:out_buffer <= mem22[12];
				13:out_buffer <= mem22[13];
				14:out_buffer <= mem22[14];
				15:out_buffer <= mem22[15];
				16:out_buffer <= mem22[16];
				17:out_buffer <= mem22[17];
				18:out_buffer <= mem22[18];
				19:out_buffer <= mem22[19];
				20:out_buffer <= mem22[20];
				21:out_buffer <= mem22[21];
				22:out_buffer <= mem22[22];
				23:out_buffer <= mem22[23];
				24:out_buffer <= mem22[24];
				25:out_buffer <= mem22[25];
				26:out_buffer <= mem22[26];
				27:out_buffer <= mem22[27];
				28:out_buffer <= mem22[28];
				29:out_buffer <= mem22[29];
			endcase
			
			23:
			case(addr)
				0:out_buffer <= mem23[0];
				1:out_buffer <= mem23[1];
				2:out_buffer <= mem23[2];
				3:out_buffer <= mem23[3];
				4:out_buffer <= mem23[4];
				5:out_buffer <= mem23[5];
				6:out_buffer <= mem23[6];
				7:out_buffer <= mem23[7];
				8:out_buffer <= mem23[8];
				9:out_buffer <= mem23[9];
				10:out_buffer <= mem23[10];
				11:out_buffer <= mem23[11];
				12:out_buffer <= mem23[12];
				13:out_buffer <= mem23[13];
				14:out_buffer <= mem23[14];
				15:out_buffer <= mem23[15];
				16:out_buffer <= mem23[16];
				17:out_buffer <= mem23[17];
				18:out_buffer <= mem23[18];
				19:out_buffer <= mem23[19];
				20:out_buffer <= mem23[20];
				21:out_buffer <= mem23[21];
				22:out_buffer <= mem23[22];
				23:out_buffer <= mem23[23];
				24:out_buffer <= mem23[24];
				25:out_buffer <= mem23[25];
				26:out_buffer <= mem23[26];
				27:out_buffer <= mem23[27];
				28:out_buffer <= mem23[28];
				29:out_buffer <= mem23[29];
			endcase
			
			24:
			case(addr)
				0:out_buffer <= mem24[0];
				1:out_buffer <= mem24[1];
				2:out_buffer <= mem24[2];
				3:out_buffer <= mem24[3];
				4:out_buffer <= mem24[4];
				5:out_buffer <= mem24[5];
				6:out_buffer <= mem24[6];
				7:out_buffer <= mem24[7];
				8:out_buffer <= mem24[8];
				9:out_buffer <= mem24[9];
				10:out_buffer <= mem24[10];
				11:out_buffer <= mem24[11];
				12:out_buffer <= mem24[12];
				13:out_buffer <= mem24[13];
				14:out_buffer <= mem24[14];
				15:out_buffer <= mem24[15];
				16:out_buffer <= mem24[16];
				17:out_buffer <= mem24[17];
				18:out_buffer <= mem24[18];
				19:out_buffer <= mem24[19];
				20:out_buffer <= mem24[20];
				21:out_buffer <= mem24[21];
				22:out_buffer <= mem24[22];
				23:out_buffer <= mem24[23];
				24:out_buffer <= mem24[24];
				25:out_buffer <= mem24[25];
				26:out_buffer <= mem24[26];
				27:out_buffer <= mem24[27];
				28:out_buffer <= mem24[28];
				29:out_buffer <= mem24[29];
			endcase

			25:
			case(addr)
				0:out_buffer <= mem25[0];
				1:out_buffer <= mem25[1];
				2:out_buffer <= mem25[2];
				3:out_buffer <= mem25[3];
				4:out_buffer <= mem25[4];
				5:out_buffer <= mem25[5];
				6:out_buffer <= mem25[6];
				7:out_buffer <= mem25[7];
				8:out_buffer <= mem25[8];
				9:out_buffer <= mem25[9];
				10:out_buffer <= mem25[10];
				11:out_buffer <= mem25[11];
				12:out_buffer <= mem25[12];
				13:out_buffer <= mem25[13];
				14:out_buffer <= mem25[14];
				15:out_buffer <= mem25[15];
				16:out_buffer <= mem25[16];
				17:out_buffer <= mem25[17];
				18:out_buffer <= mem25[18];
				19:out_buffer <= mem25[19];
				20:out_buffer <= mem25[20];
				21:out_buffer <= mem25[21];
				22:out_buffer <= mem25[22];
				23:out_buffer <= mem25[23];
				24:out_buffer <= mem25[24];
				25:out_buffer <= mem25[25];
				26:out_buffer <= mem25[26];
				27:out_buffer <= mem25[27];
				28:out_buffer <= mem25[28];
				29:out_buffer <= mem25[29];
			endcase
			
			26:
			case(addr)
				0:out_buffer <= mem26[0];
				1:out_buffer <= mem26[1];
				2:out_buffer <= mem26[2];
				3:out_buffer <= mem26[3];
				4:out_buffer <= mem26[4];
				5:out_buffer <= mem26[5];
				6:out_buffer <= mem26[6];
				7:out_buffer <= mem26[7];
				8:out_buffer <= mem26[8];
				9:out_buffer <= mem26[9];
				10:out_buffer <= mem26[10];
				11:out_buffer <= mem26[11];
				12:out_buffer <= mem26[12];
				13:out_buffer <= mem26[13];
				14:out_buffer <= mem26[14];
				15:out_buffer <= mem26[15];
				16:out_buffer <= mem26[16];
				17:out_buffer <= mem26[17];
				18:out_buffer <= mem26[18];
				19:out_buffer <= mem26[19];
				20:out_buffer <= mem26[20];
				21:out_buffer <= mem26[21];
				22:out_buffer <= mem26[22];
				23:out_buffer <= mem26[23];
				24:out_buffer <= mem26[24];
				25:out_buffer <= mem26[25];
				26:out_buffer <= mem26[26];
				27:out_buffer <= mem26[27];
				28:out_buffer <= mem26[28];
				29:out_buffer <= mem26[29];
			endcase

			27:
			case(addr)
				0:out_buffer <= mem27[0];
				1:out_buffer <= mem27[1];
				2:out_buffer <= mem27[2];
				3:out_buffer <= mem27[3];
				4:out_buffer <= mem27[4];
				5:out_buffer <= mem27[5];
				6:out_buffer <= mem27[6];
				7:out_buffer <= mem27[7];
				8:out_buffer <= mem27[8];
				9:out_buffer <= mem27[9];
				10:out_buffer <= mem27[10];
				11:out_buffer <= mem27[11];
				12:out_buffer <= mem27[12];
				13:out_buffer <= mem27[13];
				14:out_buffer <= mem27[14];
				15:out_buffer <= mem27[15];
				16:out_buffer <= mem27[16];
				17:out_buffer <= mem27[17];
				18:out_buffer <= mem27[18];
				19:out_buffer <= mem27[19];
				20:out_buffer <= mem27[20];
				21:out_buffer <= mem27[21];
				22:out_buffer <= mem27[22];
				23:out_buffer <= mem27[23];
				24:out_buffer <= mem27[24];
				25:out_buffer <= mem27[25];
				26:out_buffer <= mem27[26];
				27:out_buffer <= mem27[27];
				28:out_buffer <= mem27[28];
				29:out_buffer <= mem27[29];
			endcase

			28:
			case(addr)
				0:out_buffer <= mem28[0];
				1:out_buffer <= mem28[1];
				2:out_buffer <= mem28[2];
				3:out_buffer <= mem28[3];
				4:out_buffer <= mem28[4];
				5:out_buffer <= mem28[5];
				6:out_buffer <= mem28[6];
				7:out_buffer <= mem28[7];
				8:out_buffer <= mem28[8];
				9:out_buffer <= mem28[9];
				10:out_buffer <= mem28[10];
				11:out_buffer <= mem28[11];
				12:out_buffer <= mem28[12];
				13:out_buffer <= mem28[13];
				14:out_buffer <= mem28[14];
				15:out_buffer <= mem28[15];
				16:out_buffer <= mem28[16];
				17:out_buffer <= mem28[17];
				18:out_buffer <= mem28[18];
				19:out_buffer <= mem28[19];
				20:out_buffer <= mem28[20];
				21:out_buffer <= mem28[21];
				22:out_buffer <= mem28[22];
				23:out_buffer <= mem28[23];
				24:out_buffer <= mem28[24];
				25:out_buffer <= mem28[25];
				26:out_buffer <= mem28[26];
				27:out_buffer <= mem28[27];
				28:out_buffer <= mem28[28];
				29:out_buffer <= mem28[29];
			endcase

			29:
			case(addr)
				0:out_buffer <= mem29[0];
				1:out_buffer <= mem29[1];
				2:out_buffer <= mem29[2];
				3:out_buffer <= mem29[3];
				4:out_buffer <= mem29[4];
				5:out_buffer <= mem29[5];
				6:out_buffer <= mem29[6];
				7:out_buffer <= mem29[7];
				8:out_buffer <= mem29[8];
				9:out_buffer <= mem29[9];
				10:out_buffer <= mem29[10];
				11:out_buffer <= mem29[11];
				12:out_buffer <= mem29[12];
				13:out_buffer <= mem29[13];
				14:out_buffer <= mem29[14];
				15:out_buffer <= mem29[15];
				16:out_buffer <= mem29[16];
				17:out_buffer <= mem29[17];
				18:out_buffer <= mem29[18];
				19:out_buffer <= mem29[19];
				20:out_buffer <= mem29[20];
				21:out_buffer <= mem29[21];
				22:out_buffer <= mem29[22];
				23:out_buffer <= mem29[23];
				24:out_buffer <= mem29[24];
				25:out_buffer <= mem29[25];
				26:out_buffer <= mem29[26];
				27:out_buffer <= mem29[27];
				28:out_buffer <= mem29[28];
				29:out_buffer <= mem29[29];
			endcase
        endcase
    else if(wr_en)
		case (target_line)
			0:
			case(addr)
				0:mem00[0] <= data_in;
				1:mem00[1] <= data_in;
				2:mem00[2] <= data_in;
				3:mem00[3] <= data_in;
				4:mem00[4] <= data_in;
				5:mem00[5] <= data_in;
				6:mem00[6] <= data_in;
				7:mem00[7] <= data_in;
				8:mem00[8] <= data_in;
				9:mem00[9] <= data_in;
				10:mem00[10] <= data_in;
				11:mem00[11] <= data_in;
				12:mem00[12] <= data_in;
				13:mem00[13] <= data_in;
				14:mem00[14] <= data_in;
				15:mem00[15] <= data_in;
				16:mem00[16] <= data_in;
				17:mem00[17] <= data_in;
				18:mem00[18] <= data_in;
				19:mem00[19] <= data_in;
				20:mem00[20] <= data_in;
				21:mem00[21] <= data_in;
				22:mem00[22] <= data_in;
				23:mem00[23] <= data_in;
				24:mem00[24] <= data_in;
				25:mem00[25] <= data_in;
				26:mem00[26] <= data_in;
				27:mem00[27] <= data_in;
				28:mem00[28] <= data_in;
				29:mem00[29] <= data_in;
			endcase

			1:
			case(addr)
				0:mem01[0] <= data_in;
				1:mem01[1] <= data_in;
				2:mem01[2] <= data_in;
				3:mem01[3] <= data_in;
				4:mem01[4] <= data_in;
				5:mem01[5] <= data_in;
				6:mem01[6] <= data_in;
				7:mem01[7] <= data_in;
				8:mem01[8] <= data_in;
				9:mem01[9] <= data_in;
				10:mem01[10] <= data_in;
				11:mem01[11] <= data_in;
				12:mem01[12] <= data_in;
				13:mem01[13] <= data_in;
				14:mem01[14] <= data_in;
				15:mem01[15] <= data_in;
				16:mem01[16] <= data_in;
				17:mem01[17] <= data_in;
				18:mem01[18] <= data_in;
				19:mem01[19] <= data_in;
				20:mem01[20] <= data_in;
				21:mem01[21] <= data_in;
				22:mem01[22] <= data_in;
				23:mem01[23] <= data_in;
				24:mem01[24] <= data_in;
				25:mem01[25] <= data_in;
				26:mem01[26] <= data_in;
				27:mem01[27] <= data_in;
				28:mem01[28] <= data_in;
				29:mem01[29] <= data_in;
			endcase

			2:
			case(addr)
				0:mem02[0] <= data_in;
				1:mem02[1] <= data_in;
				2:mem02[2] <= data_in;
				3:mem02[3] <= data_in;
				4:mem02[4] <= data_in;
				5:mem02[5] <= data_in;
				6:mem02[6] <= data_in;
				7:mem02[7] <= data_in;
				8:mem02[8] <= data_in;
				9:mem02[9] <= data_in;
				10:mem02[10] <= data_in;
				11:mem02[11] <= data_in;
				12:mem02[12] <= data_in;
				13:mem02[13] <= data_in;
				14:mem02[14] <= data_in;
				15:mem02[15] <= data_in;
				16:mem02[16] <= data_in;
				17:mem02[17] <= data_in;
				18:mem02[18] <= data_in;
				19:mem02[19] <= data_in;
				20:mem02[20] <= data_in;
				21:mem02[21] <= data_in;
				22:mem02[22] <= data_in;
				23:mem02[23] <= data_in;
				24:mem02[24] <= data_in;
				25:mem02[25] <= data_in;
				26:mem02[26] <= data_in;
				27:mem02[27] <= data_in;
				28:mem02[28] <= data_in;
				29:mem02[29] <= data_in;
			endcase

			3:
			case(addr)
				0:mem03[0] <= data_in;
				1:mem03[1] <= data_in;
				2:mem03[2] <= data_in;
				3:mem03[3] <= data_in;
				4:mem03[4] <= data_in;
				5:mem03[5] <= data_in;
				6:mem03[6] <= data_in;
				7:mem03[7] <= data_in;
				8:mem03[8] <= data_in;
				9:mem03[9] <= data_in;
				10:mem03[10] <= data_in;
				11:mem03[11] <= data_in;
				12:mem03[12] <= data_in;
				13:mem03[13] <= data_in;
				14:mem03[14] <= data_in;
				15:mem03[15] <= data_in;
				16:mem03[16] <= data_in;
				17:mem03[17] <= data_in;
				18:mem03[18] <= data_in;
				19:mem03[19] <= data_in;
				20:mem03[20] <= data_in;
				21:mem03[21] <= data_in;
				22:mem03[22] <= data_in;
				23:mem03[23] <= data_in;
				24:mem03[24] <= data_in;
				25:mem03[25] <= data_in;
				26:mem03[26] <= data_in;
				27:mem03[27] <= data_in;
				28:mem03[28] <= data_in;
				29:mem03[29] <= data_in;
			endcase

			4:
			case(addr)
				0:mem04[0] <= data_in;
				1:mem04[1] <= data_in;
				2:mem04[2] <= data_in;
				3:mem04[3] <= data_in;
				4:mem04[4] <= data_in;
				5:mem04[5] <= data_in;
				6:mem04[6] <= data_in;
				7:mem04[7] <= data_in;
				8:mem04[8] <= data_in;
				9:mem04[9] <= data_in;
				10:mem04[10] <= data_in;
				11:mem04[11] <= data_in;
				12:mem04[12] <= data_in;
				13:mem04[13] <= data_in;
				14:mem04[14] <= data_in;
				15:mem04[15] <= data_in;
				16:mem04[16] <= data_in;
				17:mem04[17] <= data_in;
				18:mem04[18] <= data_in;
				19:mem04[19] <= data_in;
				20:mem04[20] <= data_in;
				21:mem04[21] <= data_in;
				22:mem04[22] <= data_in;
				23:mem04[23] <= data_in;
				24:mem04[24] <= data_in;
				25:mem04[25] <= data_in;
				26:mem04[26] <= data_in;
				27:mem04[27] <= data_in;
				28:mem04[28] <= data_in;
				29:mem04[29] <= data_in;
			endcase

			5:
			case(addr)
				0:mem05[0] <= data_in;
				1:mem05[1] <= data_in;
				2:mem05[2] <= data_in;
				3:mem05[3] <= data_in;
				4:mem05[4] <= data_in;
				5:mem05[5] <= data_in;
				6:mem05[6] <= data_in;
				7:mem05[7] <= data_in;
				8:mem05[8] <= data_in;
				9:mem05[9] <= data_in;
				10:mem05[10] <= data_in;
				11:mem05[11] <= data_in;
				12:mem05[12] <= data_in;
				13:mem05[13] <= data_in;
				14:mem05[14] <= data_in;
				15:mem05[15] <= data_in;
				16:mem05[16] <= data_in;
				17:mem05[17] <= data_in;
				18:mem05[18] <= data_in;
				19:mem05[19] <= data_in;
				20:mem05[20] <= data_in;
				21:mem05[21] <= data_in;
				22:mem05[22] <= data_in;
				23:mem05[23] <= data_in;
				24:mem05[24] <= data_in;
				25:mem05[25] <= data_in;
				26:mem05[26] <= data_in;
				27:mem05[27] <= data_in;
				28:mem05[28] <= data_in;
				29:mem05[29] <= data_in;
			endcase

			6:
			case(addr)
				0:mem06[0] <= data_in;
				1:mem06[1] <= data_in;
				2:mem06[2] <= data_in;
				3:mem06[3] <= data_in;
				4:mem06[4] <= data_in;
				5:mem06[5] <= data_in;
				6:mem06[6] <= data_in;
				7:mem06[7] <= data_in;
				8:mem06[8] <= data_in;
				9:mem06[9] <= data_in;
				10:mem06[10] <= data_in;
				11:mem06[11] <= data_in;
				12:mem06[12] <= data_in;
				13:mem06[13] <= data_in;
				14:mem06[14] <= data_in;
				15:mem06[15] <= data_in;
				16:mem06[16] <= data_in;
				17:mem06[17] <= data_in;
				18:mem06[18] <= data_in;
				19:mem06[19] <= data_in;
				20:mem06[20] <= data_in;
				21:mem06[21] <= data_in;
				22:mem06[22] <= data_in;
				23:mem06[23] <= data_in;
				24:mem06[24] <= data_in;
				25:mem06[25] <= data_in;
				26:mem06[26] <= data_in;
				27:mem06[27] <= data_in;
				28:mem06[28] <= data_in;
				29:mem06[29] <= data_in;
			endcase

			7:
			case(addr)
				0:mem07[0] <= data_in;
				1:mem07[1] <= data_in;
				2:mem07[2] <= data_in;
				3:mem07[3] <= data_in;
				4:mem07[4] <= data_in;
				5:mem07[5] <= data_in;
				6:mem07[6] <= data_in;
				7:mem07[7] <= data_in;
				8:mem07[8] <= data_in;
				9:mem07[9] <= data_in;
				10:mem07[10] <= data_in;
				11:mem07[11] <= data_in;
				12:mem07[12] <= data_in;
				13:mem07[13] <= data_in;
				14:mem07[14] <= data_in;
				15:mem07[15] <= data_in;
				16:mem07[16] <= data_in;
				17:mem07[17] <= data_in;
				18:mem07[18] <= data_in;
				19:mem07[19] <= data_in;
				20:mem07[20] <= data_in;
				21:mem07[21] <= data_in;
				22:mem07[22] <= data_in;
				23:mem07[23] <= data_in;
				24:mem07[24] <= data_in;
				25:mem07[25] <= data_in;
				26:mem07[26] <= data_in;
				27:mem07[27] <= data_in;
				28:mem07[28] <= data_in;
				29:mem07[29] <= data_in;
			endcase

			8:
			case(addr)
				0:mem08[0] <= data_in;
				1:mem08[1] <= data_in;
				2:mem08[2] <= data_in;
				3:mem08[3] <= data_in;
				4:mem08[4] <= data_in;
				5:mem08[5] <= data_in;
				6:mem08[6] <= data_in;
				7:mem08[7] <= data_in;
				8:mem08[8] <= data_in;
				9:mem08[9] <= data_in;
				10:mem08[10] <= data_in;
				11:mem08[11] <= data_in;
				12:mem08[12] <= data_in;
				13:mem08[13] <= data_in;
				14:mem08[14] <= data_in;
				15:mem08[15] <= data_in;
				16:mem08[16] <= data_in;
				17:mem08[17] <= data_in;
				18:mem08[18] <= data_in;
				19:mem08[19] <= data_in;
				20:mem08[20] <= data_in;
				21:mem08[21] <= data_in;
				22:mem08[22] <= data_in;
				23:mem08[23] <= data_in;
				24:mem08[24] <= data_in;
				25:mem08[25] <= data_in;
				26:mem08[26] <= data_in;
				27:mem08[27] <= data_in;
				28:mem08[28] <= data_in;
				29:mem08[29] <= data_in;
			endcase

			9:
			case(addr)
				0:mem09[0] <= data_in;
				1:mem09[1] <= data_in;
				2:mem09[2] <= data_in;
				3:mem09[3] <= data_in;
				4:mem09[4] <= data_in;
				5:mem09[5] <= data_in;
				6:mem09[6] <= data_in;
				7:mem09[7] <= data_in;
				8:mem09[8] <= data_in;
				9:mem09[9] <= data_in;
				10:mem09[10] <= data_in;
				11:mem09[11] <= data_in;
				12:mem09[12] <= data_in;
				13:mem09[13] <= data_in;
				14:mem09[14] <= data_in;
				15:mem09[15] <= data_in;
				16:mem09[16] <= data_in;
				17:mem09[17] <= data_in;
				18:mem09[18] <= data_in;
				19:mem09[19] <= data_in;
				20:mem09[20] <= data_in;
				21:mem09[21] <= data_in;
				22:mem09[22] <= data_in;
				23:mem09[23] <= data_in;
				24:mem09[24] <= data_in;
				25:mem09[25] <= data_in;
				26:mem09[26] <= data_in;
				27:mem09[27] <= data_in;
				28:mem09[28] <= data_in;
				29:mem09[29] <= data_in;
			endcase

			10:
			case(addr)
				0:mem10[0] <= data_in;
				1:mem10[1] <= data_in;
				2:mem10[2] <= data_in;
				3:mem10[3] <= data_in;
				4:mem10[4] <= data_in;
				5:mem10[5] <= data_in;
				6:mem10[6] <= data_in;
				7:mem10[7] <= data_in;
				8:mem10[8] <= data_in;
				9:mem10[9] <= data_in;
				10:mem10[10] <= data_in;
				11:mem10[11] <= data_in;
				12:mem10[12] <= data_in;
				13:mem10[13] <= data_in;
				14:mem10[14] <= data_in;
				15:mem10[15] <= data_in;
				16:mem10[16] <= data_in;
				17:mem10[17] <= data_in;
				18:mem10[18] <= data_in;
				19:mem10[19] <= data_in;
				20:mem10[20] <= data_in;
				21:mem10[21] <= data_in;
				22:mem10[22] <= data_in;
				23:mem10[23] <= data_in;
				24:mem10[24] <= data_in;
				25:mem10[25] <= data_in;
				26:mem10[26] <= data_in;
				27:mem10[27] <= data_in;
				28:mem10[28] <= data_in;
				29:mem10[29] <= data_in;
			endcase

			11:
			case(addr)
				0:mem11[0] <= data_in;
				1:mem11[1] <= data_in;
				2:mem11[2] <= data_in;
				3:mem11[3] <= data_in;
				4:mem11[4] <= data_in;
				5:mem11[5] <= data_in;
				6:mem11[6] <= data_in;
				7:mem11[7] <= data_in;
				8:mem11[8] <= data_in;
				9:mem11[9] <= data_in;
				10:mem11[10] <= data_in;
				11:mem11[11] <= data_in;
				12:mem11[12] <= data_in;
				13:mem11[13] <= data_in;
				14:mem11[14] <= data_in;
				15:mem11[15] <= data_in;
				16:mem11[16] <= data_in;
				17:mem11[17] <= data_in;
				18:mem11[18] <= data_in;
				19:mem11[19] <= data_in;
				20:mem11[20] <= data_in;
				21:mem11[21] <= data_in;
				22:mem11[22] <= data_in;
				23:mem11[23] <= data_in;
				24:mem11[24] <= data_in;
				25:mem11[25] <= data_in;
				26:mem11[26] <= data_in;
				27:mem11[27] <= data_in;
				28:mem11[28] <= data_in;
				29:mem11[29] <= data_in;
			endcase

			12:
			case(addr)
				0:mem12[0] <= data_in;
				1:mem12[1] <= data_in;
				2:mem12[2] <= data_in;
				3:mem12[3] <= data_in;
				4:mem12[4] <= data_in;
				5:mem12[5] <= data_in;
				6:mem12[6] <= data_in;
				7:mem12[7] <= data_in;
				8:mem12[8] <= data_in;
				9:mem12[9] <= data_in;
				10:mem12[10] <= data_in;
				11:mem12[11] <= data_in;
				12:mem12[12] <= data_in;
				13:mem12[13] <= data_in;
				14:mem12[14] <= data_in;
				15:mem12[15] <= data_in;
				16:mem12[16] <= data_in;
				17:mem12[17] <= data_in;
				18:mem12[18] <= data_in;
				19:mem12[19] <= data_in;
				20:mem12[20] <= data_in;
				21:mem12[21] <= data_in;
				22:mem12[22] <= data_in;
				23:mem12[23] <= data_in;
				24:mem12[24] <= data_in;
				25:mem12[25] <= data_in;
				26:mem12[26] <= data_in;
				27:mem12[27] <= data_in;
				28:mem12[28] <= data_in;
				29:mem12[29] <= data_in;
			endcase

			13:
			case(addr)
				0:mem13[0] <= data_in;
				1:mem13[1] <= data_in;
				2:mem13[2] <= data_in;
				3:mem13[3] <= data_in;
				4:mem13[4] <= data_in;
				5:mem13[5] <= data_in;
				6:mem13[6] <= data_in;
				7:mem13[7] <= data_in;
				8:mem13[8] <= data_in;
				9:mem13[9] <= data_in;
				10:mem13[10] <= data_in;
				11:mem13[11] <= data_in;
				12:mem13[12] <= data_in;
				13:mem13[13] <= data_in;
				14:mem13[14] <= data_in;
				15:mem13[15] <= data_in;
				16:mem13[16] <= data_in;
				17:mem13[17] <= data_in;
				18:mem13[18] <= data_in;
				19:mem13[19] <= data_in;
				20:mem13[20] <= data_in;
				21:mem13[21] <= data_in;
				22:mem13[22] <= data_in;
				23:mem13[23] <= data_in;
				24:mem13[24] <= data_in;
				25:mem13[25] <= data_in;
				26:mem13[26] <= data_in;
				27:mem13[27] <= data_in;
				28:mem13[28] <= data_in;
				29:mem13[29] <= data_in;
			endcase

			14:
			case(addr)
				0:mem14[0] <= data_in;
				1:mem14[1] <= data_in;
				2:mem14[2] <= data_in;
				3:mem14[3] <= data_in;
				4:mem14[4] <= data_in;
				5:mem14[5] <= data_in;
				6:mem14[6] <= data_in;
				7:mem14[7] <= data_in;
				8:mem14[8] <= data_in;
				9:mem14[9] <= data_in;
				10:mem14[10] <= data_in;
				11:mem14[11] <= data_in;
				12:mem14[12] <= data_in;
				13:mem14[13] <= data_in;
				14:mem14[14] <= data_in;
				15:mem14[15] <= data_in;
				16:mem14[16] <= data_in;
				17:mem14[17] <= data_in;
				18:mem14[18] <= data_in;
				19:mem14[19] <= data_in;
				20:mem14[20] <= data_in;
				21:mem14[21] <= data_in;
				22:mem14[22] <= data_in;
				23:mem14[23] <= data_in;
				24:mem14[24] <= data_in;
				25:mem14[25] <= data_in;
				26:mem14[26] <= data_in;
				27:mem14[27] <= data_in;
				28:mem14[28] <= data_in;
				29:mem14[29] <= data_in;
			endcase

			15:
			case(addr)
				0:mem15[0] <= data_in;
				1:mem15[1] <= data_in;
				2:mem15[2] <= data_in;
				3:mem15[3] <= data_in;
				4:mem15[4] <= data_in;
				5:mem15[5] <= data_in;
				6:mem15[6] <= data_in;
				7:mem15[7] <= data_in;
				8:mem15[8] <= data_in;
				9:mem15[9] <= data_in;
				10:mem15[10] <= data_in;
				11:mem15[11] <= data_in;
				12:mem15[12] <= data_in;
				13:mem15[13] <= data_in;
				14:mem15[14] <= data_in;
				15:mem15[15] <= data_in;
				16:mem15[16] <= data_in;
				17:mem15[17] <= data_in;
				18:mem15[18] <= data_in;
				19:mem15[19] <= data_in;
				20:mem15[20] <= data_in;
				21:mem15[21] <= data_in;
				22:mem15[22] <= data_in;
				23:mem15[23] <= data_in;
				24:mem15[24] <= data_in;
				25:mem15[25] <= data_in;
				26:mem15[26] <= data_in;
				27:mem15[27] <= data_in;
				28:mem15[28] <= data_in;
				29:mem15[29] <= data_in;
			endcase

			16:
			case(addr)
				0:mem16[0] <= data_in;
				1:mem16[1] <= data_in;
				2:mem16[2] <= data_in;
				3:mem16[3] <= data_in;
				4:mem16[4] <= data_in;
				5:mem16[5] <= data_in;
				6:mem16[6] <= data_in;
				7:mem16[7] <= data_in;
				8:mem16[8] <= data_in;
				9:mem16[9] <= data_in;
				10:mem16[10] <= data_in;
				11:mem16[11] <= data_in;
				12:mem16[12] <= data_in;
				13:mem16[13] <= data_in;
				14:mem16[14] <= data_in;
				15:mem16[15] <= data_in;
				16:mem16[16] <= data_in;
				17:mem16[17] <= data_in;
				18:mem16[18] <= data_in;
				19:mem16[19] <= data_in;
				20:mem16[20] <= data_in;
				21:mem16[21] <= data_in;
				22:mem16[22] <= data_in;
				23:mem16[23] <= data_in;
				24:mem16[24] <= data_in;
				25:mem16[25] <= data_in;
				26:mem16[26] <= data_in;
				27:mem16[27] <= data_in;
				28:mem16[28] <= data_in;
				29:mem16[29] <= data_in;
			endcase

			17:
			case(addr)
				0:mem17[0] <= data_in;
				1:mem17[1] <= data_in;
				2:mem17[2] <= data_in;
				3:mem17[3] <= data_in;
				4:mem17[4] <= data_in;
				5:mem17[5] <= data_in;
				6:mem17[6] <= data_in;
				7:mem17[7] <= data_in;
				8:mem17[8] <= data_in;
				9:mem17[9] <= data_in;
				10:mem17[10] <= data_in;
				11:mem17[11] <= data_in;
				12:mem17[12] <= data_in;
				13:mem17[13] <= data_in;
				14:mem17[14] <= data_in;
				15:mem17[15] <= data_in;
				16:mem17[16] <= data_in;
				17:mem17[17] <= data_in;
				18:mem17[18] <= data_in;
				19:mem17[19] <= data_in;
				20:mem17[20] <= data_in;
				21:mem17[21] <= data_in;
				22:mem17[22] <= data_in;
				23:mem17[23] <= data_in;
				24:mem17[24] <= data_in;
				25:mem17[25] <= data_in;
				26:mem17[26] <= data_in;
				27:mem17[27] <= data_in;
				28:mem17[28] <= data_in;
				29:mem17[29] <= data_in;
			endcase

			18:
			case(addr)
				0:mem18[0] <= data_in;
				1:mem18[1] <= data_in;
				2:mem18[2] <= data_in;
				3:mem18[3] <= data_in;
				4:mem18[4] <= data_in;
				5:mem18[5] <= data_in;
				6:mem18[6] <= data_in;
				7:mem18[7] <= data_in;
				8:mem18[8] <= data_in;
				9:mem18[9] <= data_in;
				10:mem18[10] <= data_in;
				11:mem18[11] <= data_in;
				12:mem18[12] <= data_in;
				13:mem18[13] <= data_in;
				14:mem18[14] <= data_in;
				15:mem18[15] <= data_in;
				16:mem18[16] <= data_in;
				17:mem18[17] <= data_in;
				18:mem18[18] <= data_in;
				19:mem18[19] <= data_in;
				20:mem18[20] <= data_in;
				21:mem18[21] <= data_in;
				22:mem18[22] <= data_in;
				23:mem18[23] <= data_in;
				24:mem18[24] <= data_in;
				25:mem18[25] <= data_in;
				26:mem18[26] <= data_in;
				27:mem18[27] <= data_in;
				28:mem18[28] <= data_in;
				29:mem18[29] <= data_in;
			endcase

			19:
			case(addr)
				0:mem19[0] <= data_in;
				1:mem19[1] <= data_in;
				2:mem19[2] <= data_in;
				3:mem19[3] <= data_in;
				4:mem19[4] <= data_in;
				5:mem19[5] <= data_in;
				6:mem19[6] <= data_in;
				7:mem19[7] <= data_in;
				8:mem19[8] <= data_in;
				9:mem19[9] <= data_in;
				10:mem19[10] <= data_in;
				11:mem19[11] <= data_in;
				12:mem19[12] <= data_in;
				13:mem19[13] <= data_in;
				14:mem19[14] <= data_in;
				15:mem19[15] <= data_in;
				16:mem19[16] <= data_in;
				17:mem19[17] <= data_in;
				18:mem19[18] <= data_in;
				19:mem19[19] <= data_in;
				20:mem19[20] <= data_in;
				21:mem19[21] <= data_in;
				22:mem19[22] <= data_in;
				23:mem19[23] <= data_in;
				24:mem19[24] <= data_in;
				25:mem19[25] <= data_in;
				26:mem19[26] <= data_in;
				27:mem19[27] <= data_in;
				28:mem19[28] <= data_in;
				29:mem19[29] <= data_in;
			endcase

			20:
			case(addr)
				0:mem20[0] <= data_in;
				1:mem20[1] <= data_in;
				2:mem20[2] <= data_in;
				3:mem20[3] <= data_in;
				4:mem20[4] <= data_in;
				5:mem20[5] <= data_in;
				6:mem20[6] <= data_in;
				7:mem20[7] <= data_in;
				8:mem20[8] <= data_in;
				9:mem20[9] <= data_in;
				10:mem20[10] <= data_in;
				11:mem20[11] <= data_in;
				12:mem20[12] <= data_in;
				13:mem20[13] <= data_in;
				14:mem20[14] <= data_in;
				15:mem20[15] <= data_in;
				16:mem20[16] <= data_in;
				17:mem20[17] <= data_in;
				18:mem20[18] <= data_in;
				19:mem20[19] <= data_in;
				20:mem20[20] <= data_in;
				21:mem20[21] <= data_in;
				22:mem20[22] <= data_in;
				23:mem20[23] <= data_in;
				24:mem20[24] <= data_in;
				25:mem20[25] <= data_in;
				26:mem20[26] <= data_in;
				27:mem20[27] <= data_in;
				28:mem20[28] <= data_in;
				29:mem20[29] <= data_in;
			endcase

			21:
			case(addr)
				0:mem21[0] <= data_in;
				1:mem21[1] <= data_in;
				2:mem21[2] <= data_in;
				3:mem21[3] <= data_in;
				4:mem21[4] <= data_in;
				5:mem21[5] <= data_in;
				6:mem21[6] <= data_in;
				7:mem21[7] <= data_in;
				8:mem21[8] <= data_in;
				9:mem21[9] <= data_in;
				10:mem21[10] <= data_in;
				11:mem21[11] <= data_in;
				12:mem21[12] <= data_in;
				13:mem21[13] <= data_in;
				14:mem21[14] <= data_in;
				15:mem21[15] <= data_in;
				16:mem21[16] <= data_in;
				17:mem21[17] <= data_in;
				18:mem21[18] <= data_in;
				19:mem21[19] <= data_in;
				20:mem21[20] <= data_in;
				21:mem21[21] <= data_in;
				22:mem21[22] <= data_in;
				23:mem21[23] <= data_in;
				24:mem21[24] <= data_in;
				25:mem21[25] <= data_in;
				26:mem21[26] <= data_in;
				27:mem21[27] <= data_in;
				28:mem21[28] <= data_in;
				29:mem21[29] <= data_in;
			endcase

			22:
			case(addr)
				0:mem22[0] <= data_in;
				1:mem22[1] <= data_in;
				2:mem22[2] <= data_in;
				3:mem22[3] <= data_in;
				4:mem22[4] <= data_in;
				5:mem22[5] <= data_in;
				6:mem22[6] <= data_in;
				7:mem22[7] <= data_in;
				8:mem22[8] <= data_in;
				9:mem22[9] <= data_in;
				10:mem22[10] <= data_in;
				11:mem22[11] <= data_in;
				12:mem22[12] <= data_in;
				13:mem22[13] <= data_in;
				14:mem22[14] <= data_in;
				15:mem22[15] <= data_in;
				16:mem22[16] <= data_in;
				17:mem22[17] <= data_in;
				18:mem22[18] <= data_in;
				19:mem22[19] <= data_in;
				20:mem22[20] <= data_in;
				21:mem22[21] <= data_in;
				22:mem22[22] <= data_in;
				23:mem22[23] <= data_in;
				24:mem22[24] <= data_in;
				25:mem22[25] <= data_in;
				26:mem22[26] <= data_in;
				27:mem22[27] <= data_in;
				28:mem22[28] <= data_in;
				29:mem22[29] <= data_in;
			endcase

			23:
			case(addr)
				0:mem23[0] <= data_in;
				1:mem23[1] <= data_in;
				2:mem23[2] <= data_in;
				3:mem23[3] <= data_in;
				4:mem23[4] <= data_in;
				5:mem23[5] <= data_in;
				6:mem23[6] <= data_in;
				7:mem23[7] <= data_in;
				8:mem23[8] <= data_in;
				9:mem23[9] <= data_in;
				10:mem23[10] <= data_in;
				11:mem23[11] <= data_in;
				12:mem23[12] <= data_in;
				13:mem23[13] <= data_in;
				14:mem23[14] <= data_in;
				15:mem23[15] <= data_in;
				16:mem23[16] <= data_in;
				17:mem23[17] <= data_in;
				18:mem23[18] <= data_in;
				19:mem23[19] <= data_in;
				20:mem23[20] <= data_in;
				21:mem23[21] <= data_in;
				22:mem23[22] <= data_in;
				23:mem23[23] <= data_in;
				24:mem23[24] <= data_in;
				25:mem23[25] <= data_in;
				26:mem23[26] <= data_in;
				27:mem23[27] <= data_in;
				28:mem23[28] <= data_in;
				29:mem23[29] <= data_in;
			endcase

			24:
			case(addr)
				0:mem24[0] <= data_in;
				1:mem24[1] <= data_in;
				2:mem24[2] <= data_in;
				3:mem24[3] <= data_in;
				4:mem24[4] <= data_in;
				5:mem24[5] <= data_in;
				6:mem24[6] <= data_in;
				7:mem24[7] <= data_in;
				8:mem24[8] <= data_in;
				9:mem24[9] <= data_in;
				10:mem24[10] <= data_in;
				11:mem24[11] <= data_in;
				12:mem24[12] <= data_in;
				13:mem24[13] <= data_in;
				14:mem24[14] <= data_in;
				15:mem24[15] <= data_in;
				16:mem24[16] <= data_in;
				17:mem24[17] <= data_in;
				18:mem24[18] <= data_in;
				19:mem24[19] <= data_in;
				20:mem24[20] <= data_in;
				21:mem24[21] <= data_in;
				22:mem24[22] <= data_in;
				23:mem24[23] <= data_in;
				24:mem24[24] <= data_in;
				25:mem24[25] <= data_in;
				26:mem24[26] <= data_in;
				27:mem24[27] <= data_in;
				28:mem24[28] <= data_in;
				29:mem24[29] <= data_in;
			endcase

			25:
			case(addr)
				0:mem25[0] <= data_in;
				1:mem25[1] <= data_in;
				2:mem25[2] <= data_in;
				3:mem25[3] <= data_in;
				4:mem25[4] <= data_in;
				5:mem25[5] <= data_in;
				6:mem25[6] <= data_in;
				7:mem25[7] <= data_in;
				8:mem25[8] <= data_in;
				9:mem25[9] <= data_in;
				10:mem25[10] <= data_in;
				11:mem25[11] <= data_in;
				12:mem25[12] <= data_in;
				13:mem25[13] <= data_in;
				14:mem25[14] <= data_in;
				15:mem25[15] <= data_in;
				16:mem25[16] <= data_in;
				17:mem25[17] <= data_in;
				18:mem25[18] <= data_in;
				19:mem25[19] <= data_in;
				20:mem25[20] <= data_in;
				21:mem25[21] <= data_in;
				22:mem25[22] <= data_in;
				23:mem25[23] <= data_in;
				24:mem25[24] <= data_in;
				25:mem25[25] <= data_in;
				26:mem25[26] <= data_in;
				27:mem25[27] <= data_in;
				28:mem25[28] <= data_in;
				29:mem25[29] <= data_in;
			endcase

			26:
			case(addr)
				0:mem26[0] <= data_in;
				1:mem26[1] <= data_in;
				2:mem26[2] <= data_in;
				3:mem26[3] <= data_in;
				4:mem26[4] <= data_in;
				5:mem26[5] <= data_in;
				6:mem26[6] <= data_in;
				7:mem26[7] <= data_in;
				8:mem26[8] <= data_in;
				9:mem26[9] <= data_in;
				10:mem26[10] <= data_in;
				11:mem26[11] <= data_in;
				12:mem26[12] <= data_in;
				13:mem26[13] <= data_in;
				14:mem26[14] <= data_in;
				15:mem26[15] <= data_in;
				16:mem26[16] <= data_in;
				17:mem26[17] <= data_in;
				18:mem26[18] <= data_in;
				19:mem26[19] <= data_in;
				20:mem26[20] <= data_in;
				21:mem26[21] <= data_in;
				22:mem26[22] <= data_in;
				23:mem26[23] <= data_in;
				24:mem26[24] <= data_in;
				25:mem26[25] <= data_in;
				26:mem26[26] <= data_in;
				27:mem26[27] <= data_in;
				28:mem26[28] <= data_in;
				29:mem26[29] <= data_in;
			endcase

			27:
			case(addr)
				0:mem27[0] <= data_in;
				1:mem27[1] <= data_in;
				2:mem27[2] <= data_in;
				3:mem27[3] <= data_in;
				4:mem27[4] <= data_in;
				5:mem27[5] <= data_in;
				6:mem27[6] <= data_in;
				7:mem27[7] <= data_in;
				8:mem27[8] <= data_in;
				9:mem27[9] <= data_in;
				10:mem27[10] <= data_in;
				11:mem27[11] <= data_in;
				12:mem27[12] <= data_in;
				13:mem27[13] <= data_in;
				14:mem27[14] <= data_in;
				15:mem27[15] <= data_in;
				16:mem27[16] <= data_in;
				17:mem27[17] <= data_in;
				18:mem27[18] <= data_in;
				19:mem27[19] <= data_in;
				20:mem27[20] <= data_in;
				21:mem27[21] <= data_in;
				22:mem27[22] <= data_in;
				23:mem27[23] <= data_in;
				24:mem27[24] <= data_in;
				25:mem27[25] <= data_in;
				26:mem27[26] <= data_in;
				27:mem27[27] <= data_in;
				28:mem27[28] <= data_in;
				29:mem27[29] <= data_in;
			endcase

			28:
			case(addr)
				0:mem28[0] <= data_in;
				1:mem28[1] <= data_in;
				2:mem28[2] <= data_in;
				3:mem28[3] <= data_in;
				4:mem28[4] <= data_in;
				5:mem28[5] <= data_in;
				6:mem28[6] <= data_in;
				7:mem28[7] <= data_in;
				8:mem28[8] <= data_in;
				9:mem28[9] <= data_in;
				10:mem28[10] <= data_in;
				11:mem28[11] <= data_in;
				12:mem28[12] <= data_in;
				13:mem28[13] <= data_in;
				14:mem28[14] <= data_in;
				15:mem28[15] <= data_in;
				16:mem28[16] <= data_in;
				17:mem28[17] <= data_in;
				18:mem28[18] <= data_in;
				19:mem28[19] <= data_in;
				20:mem28[20] <= data_in;
				21:mem28[21] <= data_in;
				22:mem28[22] <= data_in;
				23:mem28[23] <= data_in;
				24:mem28[24] <= data_in;
				25:mem28[25] <= data_in;
				26:mem28[26] <= data_in;
				27:mem28[27] <= data_in;
				28:mem28[28] <= data_in;
				29:mem28[29] <= data_in;
			endcase

			29:
			case(addr)
				0:mem29[0] <= data_in;
				1:mem29[1] <= data_in;
				2:mem29[2] <= data_in;
				3:mem29[3] <= data_in;
				4:mem29[4] <= data_in;
				5:mem29[5] <= data_in;
				6:mem29[6] <= data_in;
				7:mem29[7] <= data_in;
				8:mem29[8] <= data_in;
				9:mem29[9] <= data_in;
				10:mem29[10] <= data_in;
				11:mem29[11] <= data_in;
				12:mem29[12] <= data_in;
				13:mem29[13] <= data_in;
				14:mem29[14] <= data_in;
				15:mem29[15] <= data_in;
				16:mem29[16] <= data_in;
				17:mem29[17] <= data_in;
				18:mem29[18] <= data_in;
				19:mem29[19] <= data_in;
				20:mem29[20] <= data_in;
				21:mem29[21] <= data_in;
				22:mem29[22] <= data_in;
				23:mem29[23] <= data_in;
				24:mem29[24] <= data_in;
				25:mem29[25] <= data_in;
				26:mem29[26] <= data_in;
				27:mem29[27] <= data_in;
				28:mem29[28] <= data_in;
				29:mem29[29] <= data_in;
			endcase
            //default:
        endcase
    else
        out_buffer <= 9'bz;//读写均无效时，为高阻态。若不加此句，时序会出现问题
end

assign out = out_buffer;

endmodule