`timescale 1ns / 1ps
// max pooling

module pooling(
    input clk,
    input rst_n,
    // data
    input 

    output 
)

endmodule
